.INIT_00(INIT[  0*256 +: 256]),
.INIT_01(INIT[  1*256 +: 256]),
.INIT_02(INIT[  2*256 +: 256]),
.INIT_03(INIT[  3*256 +: 256]),
.INIT_04(INIT[  4*256 +: 256]),
.INIT_05(INIT[  5*256 +: 256]),
.INIT_06(INIT[  6*256 +: 256]),
.INIT_07(INIT[  7*256 +: 256]),
.INIT_08(INIT[  8*256 +: 256]),
.INIT_09(INIT[  9*256 +: 256]),
.INIT_0A(INIT[ 10*256 +: 256]),
.INIT_0B(INIT[ 11*256 +: 256]),
.INIT_0C(INIT[ 12*256 +: 256]),
.INIT_0D(INIT[ 13*256 +: 256]),
.INIT_0E(INIT[ 14*256 +: 256]),
.INIT_0F(INIT[ 15*256 +: 256]),
.INIT_10(INIT[ 16*256 +: 256]),
.INIT_11(INIT[ 17*256 +: 256]),
.INIT_12(INIT[ 18*256 +: 256]),
.INIT_13(INIT[ 19*256 +: 256]),
.INIT_14(INIT[ 20*256 +: 256]),
.INIT_15(INIT[ 21*256 +: 256]),
.INIT_16(INIT[ 22*256 +: 256]),
.INIT_17(INIT[ 23*256 +: 256]),
.INIT_18(INIT[ 24*256 +: 256]),
.INIT_19(INIT[ 25*256 +: 256]),
.INIT_1A(INIT[ 26*256 +: 256]),
.INIT_1B(INIT[ 27*256 +: 256]),
.INIT_1C(INIT[ 28*256 +: 256]),
.INIT_1D(INIT[ 29*256 +: 256]),
.INIT_1E(INIT[ 30*256 +: 256]),
.INIT_1F(INIT[ 31*256 +: 256]),
.INIT_20(INIT[ 32*256 +: 256]),
.INIT_21(INIT[ 33*256 +: 256]),
.INIT_22(INIT[ 34*256 +: 256]),
.INIT_23(INIT[ 35*256 +: 256]),
.INIT_24(INIT[ 36*256 +: 256]),
.INIT_25(INIT[ 37*256 +: 256]),
.INIT_26(INIT[ 38*256 +: 256]),
.INIT_27(INIT[ 39*256 +: 256]),
.INIT_28(INIT[ 40*256 +: 256]),
.INIT_29(INIT[ 41*256 +: 256]),
.INIT_2A(INIT[ 42*256 +: 256]),
.INIT_2B(INIT[ 43*256 +: 256]),
.INIT_2C(INIT[ 44*256 +: 256]),
.INIT_2D(INIT[ 45*256 +: 256]),
.INIT_2E(INIT[ 46*256 +: 256]),
.INIT_2F(INIT[ 47*256 +: 256]),
.INIT_30(INIT[ 48*256 +: 256]),
.INIT_31(INIT[ 49*256 +: 256]),
.INIT_32(INIT[ 50*256 +: 256]),
.INIT_33(INIT[ 51*256 +: 256]),
.INIT_34(INIT[ 52*256 +: 256]),
.INIT_35(INIT[ 53*256 +: 256]),
.INIT_36(INIT[ 54*256 +: 256]),
.INIT_37(INIT[ 55*256 +: 256]),
.INIT_38(INIT[ 56*256 +: 256]),
.INIT_39(INIT[ 57*256 +: 256]),
.INIT_3A(INIT[ 58*256 +: 256]),
.INIT_3B(INIT[ 59*256 +: 256]),
.INIT_3C(INIT[ 60*256 +: 256]),
.INIT_3D(INIT[ 61*256 +: 256]),
.INIT_3E(INIT[ 62*256 +: 256]),
.INIT_3F(INIT[ 63*256 +: 256]),
