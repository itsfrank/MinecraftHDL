.INITP_00({INIT[255*9+8], INIT[254*9+8], INIT[253*9+8], INIT[252*9+8], 
           INIT[251*9+8], INIT[250*9+8], INIT[249*9+8], INIT[248*9+8], 
           INIT[247*9+8], INIT[246*9+8], INIT[245*9+8], INIT[244*9+8], 
           INIT[243*9+8], INIT[242*9+8], INIT[241*9+8], INIT[240*9+8], 
           INIT[239*9+8], INIT[238*9+8], INIT[237*9+8], INIT[236*9+8], 
           INIT[235*9+8], INIT[234*9+8], INIT[233*9+8], INIT[232*9+8], 
           INIT[231*9+8], INIT[230*9+8], INIT[229*9+8], INIT[228*9+8], 
           INIT[227*9+8], INIT[226*9+8], INIT[225*9+8], INIT[224*9+8], 
           INIT[223*9+8], INIT[222*9+8], INIT[221*9+8], INIT[220*9+8], 
           INIT[219*9+8], INIT[218*9+8], INIT[217*9+8], INIT[216*9+8], 
           INIT[215*9+8], INIT[214*9+8], INIT[213*9+8], INIT[212*9+8], 
           INIT[211*9+8], INIT[210*9+8], INIT[209*9+8], INIT[208*9+8], 
           INIT[207*9+8], INIT[206*9+8], INIT[205*9+8], INIT[204*9+8], 
           INIT[203*9+8], INIT[202*9+8], INIT[201*9+8], INIT[200*9+8], 
           INIT[199*9+8], INIT[198*9+8], INIT[197*9+8], INIT[196*9+8], 
           INIT[195*9+8], INIT[194*9+8], INIT[193*9+8], INIT[192*9+8], 
           INIT[191*9+8], INIT[190*9+8], INIT[189*9+8], INIT[188*9+8], 
           INIT[187*9+8], INIT[186*9+8], INIT[185*9+8], INIT[184*9+8], 
           INIT[183*9+8], INIT[182*9+8], INIT[181*9+8], INIT[180*9+8], 
           INIT[179*9+8], INIT[178*9+8], INIT[177*9+8], INIT[176*9+8], 
           INIT[175*9+8], INIT[174*9+8], INIT[173*9+8], INIT[172*9+8], 
           INIT[171*9+8], INIT[170*9+8], INIT[169*9+8], INIT[168*9+8], 
           INIT[167*9+8], INIT[166*9+8], INIT[165*9+8], INIT[164*9+8], 
           INIT[163*9+8], INIT[162*9+8], INIT[161*9+8], INIT[160*9+8], 
           INIT[159*9+8], INIT[158*9+8], INIT[157*9+8], INIT[156*9+8], 
           INIT[155*9+8], INIT[154*9+8], INIT[153*9+8], INIT[152*9+8], 
           INIT[151*9+8], INIT[150*9+8], INIT[149*9+8], INIT[148*9+8], 
           INIT[147*9+8], INIT[146*9+8], INIT[145*9+8], INIT[144*9+8], 
           INIT[143*9+8], INIT[142*9+8], INIT[141*9+8], INIT[140*9+8], 
           INIT[139*9+8], INIT[138*9+8], INIT[137*9+8], INIT[136*9+8], 
           INIT[135*9+8], INIT[134*9+8], INIT[133*9+8], INIT[132*9+8], 
           INIT[131*9+8], INIT[130*9+8], INIT[129*9+8], INIT[128*9+8], 
           INIT[127*9+8], INIT[126*9+8], INIT[125*9+8], INIT[124*9+8], 
           INIT[123*9+8], INIT[122*9+8], INIT[121*9+8], INIT[120*9+8], 
           INIT[119*9+8], INIT[118*9+8], INIT[117*9+8], INIT[116*9+8], 
           INIT[115*9+8], INIT[114*9+8], INIT[113*9+8], INIT[112*9+8], 
           INIT[111*9+8], INIT[110*9+8], INIT[109*9+8], INIT[108*9+8], 
           INIT[107*9+8], INIT[106*9+8], INIT[105*9+8], INIT[104*9+8], 
           INIT[103*9+8], INIT[102*9+8], INIT[101*9+8], INIT[100*9+8], 
           INIT[ 99*9+8], INIT[ 98*9+8], INIT[ 97*9+8], INIT[ 96*9+8], 
           INIT[ 95*9+8], INIT[ 94*9+8], INIT[ 93*9+8], INIT[ 92*9+8], 
           INIT[ 91*9+8], INIT[ 90*9+8], INIT[ 89*9+8], INIT[ 88*9+8], 
           INIT[ 87*9+8], INIT[ 86*9+8], INIT[ 85*9+8], INIT[ 84*9+8], 
           INIT[ 83*9+8], INIT[ 82*9+8], INIT[ 81*9+8], INIT[ 80*9+8], 
           INIT[ 79*9+8], INIT[ 78*9+8], INIT[ 77*9+8], INIT[ 76*9+8], 
           INIT[ 75*9+8], INIT[ 74*9+8], INIT[ 73*9+8], INIT[ 72*9+8], 
           INIT[ 71*9+8], INIT[ 70*9+8], INIT[ 69*9+8], INIT[ 68*9+8], 
           INIT[ 67*9+8], INIT[ 66*9+8], INIT[ 65*9+8], INIT[ 64*9+8], 
           INIT[ 63*9+8], INIT[ 62*9+8], INIT[ 61*9+8], INIT[ 60*9+8], 
           INIT[ 59*9+8], INIT[ 58*9+8], INIT[ 57*9+8], INIT[ 56*9+8], 
           INIT[ 55*9+8], INIT[ 54*9+8], INIT[ 53*9+8], INIT[ 52*9+8], 
           INIT[ 51*9+8], INIT[ 50*9+8], INIT[ 49*9+8], INIT[ 48*9+8], 
           INIT[ 47*9+8], INIT[ 46*9+8], INIT[ 45*9+8], INIT[ 44*9+8], 
           INIT[ 43*9+8], INIT[ 42*9+8], INIT[ 41*9+8], INIT[ 40*9+8], 
           INIT[ 39*9+8], INIT[ 38*9+8], INIT[ 37*9+8], INIT[ 36*9+8], 
           INIT[ 35*9+8], INIT[ 34*9+8], INIT[ 33*9+8], INIT[ 32*9+8], 
           INIT[ 31*9+8], INIT[ 30*9+8], INIT[ 29*9+8], INIT[ 28*9+8], 
           INIT[ 27*9+8], INIT[ 26*9+8], INIT[ 25*9+8], INIT[ 24*9+8], 
           INIT[ 23*9+8], INIT[ 22*9+8], INIT[ 21*9+8], INIT[ 20*9+8], 
           INIT[ 19*9+8], INIT[ 18*9+8], INIT[ 17*9+8], INIT[ 16*9+8], 
           INIT[ 15*9+8], INIT[ 14*9+8], INIT[ 13*9+8], INIT[ 12*9+8], 
           INIT[ 11*9+8], INIT[ 10*9+8], INIT[  9*9+8], INIT[  8*9+8], 
           INIT[  7*9+8], INIT[  6*9+8], INIT[  5*9+8], INIT[  4*9+8], 
           INIT[  3*9+8], INIT[  2*9+8], INIT[  1*9+8], INIT[  0*9+8]}),
.INITP_01({INIT[511*9+8], INIT[510*9+8], INIT[509*9+8], INIT[508*9+8], 
           INIT[507*9+8], INIT[506*9+8], INIT[505*9+8], INIT[504*9+8], 
           INIT[503*9+8], INIT[502*9+8], INIT[501*9+8], INIT[500*9+8], 
           INIT[499*9+8], INIT[498*9+8], INIT[497*9+8], INIT[496*9+8], 
           INIT[495*9+8], INIT[494*9+8], INIT[493*9+8], INIT[492*9+8], 
           INIT[491*9+8], INIT[490*9+8], INIT[489*9+8], INIT[488*9+8], 
           INIT[487*9+8], INIT[486*9+8], INIT[485*9+8], INIT[484*9+8], 
           INIT[483*9+8], INIT[482*9+8], INIT[481*9+8], INIT[480*9+8], 
           INIT[479*9+8], INIT[478*9+8], INIT[477*9+8], INIT[476*9+8], 
           INIT[475*9+8], INIT[474*9+8], INIT[473*9+8], INIT[472*9+8], 
           INIT[471*9+8], INIT[470*9+8], INIT[469*9+8], INIT[468*9+8], 
           INIT[467*9+8], INIT[466*9+8], INIT[465*9+8], INIT[464*9+8], 
           INIT[463*9+8], INIT[462*9+8], INIT[461*9+8], INIT[460*9+8], 
           INIT[459*9+8], INIT[458*9+8], INIT[457*9+8], INIT[456*9+8], 
           INIT[455*9+8], INIT[454*9+8], INIT[453*9+8], INIT[452*9+8], 
           INIT[451*9+8], INIT[450*9+8], INIT[449*9+8], INIT[448*9+8], 
           INIT[447*9+8], INIT[446*9+8], INIT[445*9+8], INIT[444*9+8], 
           INIT[443*9+8], INIT[442*9+8], INIT[441*9+8], INIT[440*9+8], 
           INIT[439*9+8], INIT[438*9+8], INIT[437*9+8], INIT[436*9+8], 
           INIT[435*9+8], INIT[434*9+8], INIT[433*9+8], INIT[432*9+8], 
           INIT[431*9+8], INIT[430*9+8], INIT[429*9+8], INIT[428*9+8], 
           INIT[427*9+8], INIT[426*9+8], INIT[425*9+8], INIT[424*9+8], 
           INIT[423*9+8], INIT[422*9+8], INIT[421*9+8], INIT[420*9+8], 
           INIT[419*9+8], INIT[418*9+8], INIT[417*9+8], INIT[416*9+8], 
           INIT[415*9+8], INIT[414*9+8], INIT[413*9+8], INIT[412*9+8], 
           INIT[411*9+8], INIT[410*9+8], INIT[409*9+8], INIT[408*9+8], 
           INIT[407*9+8], INIT[406*9+8], INIT[405*9+8], INIT[404*9+8], 
           INIT[403*9+8], INIT[402*9+8], INIT[401*9+8], INIT[400*9+8], 
           INIT[399*9+8], INIT[398*9+8], INIT[397*9+8], INIT[396*9+8], 
           INIT[395*9+8], INIT[394*9+8], INIT[393*9+8], INIT[392*9+8], 
           INIT[391*9+8], INIT[390*9+8], INIT[389*9+8], INIT[388*9+8], 
           INIT[387*9+8], INIT[386*9+8], INIT[385*9+8], INIT[384*9+8], 
           INIT[383*9+8], INIT[382*9+8], INIT[381*9+8], INIT[380*9+8], 
           INIT[379*9+8], INIT[378*9+8], INIT[377*9+8], INIT[376*9+8], 
           INIT[375*9+8], INIT[374*9+8], INIT[373*9+8], INIT[372*9+8], 
           INIT[371*9+8], INIT[370*9+8], INIT[369*9+8], INIT[368*9+8], 
           INIT[367*9+8], INIT[366*9+8], INIT[365*9+8], INIT[364*9+8], 
           INIT[363*9+8], INIT[362*9+8], INIT[361*9+8], INIT[360*9+8], 
           INIT[359*9+8], INIT[358*9+8], INIT[357*9+8], INIT[356*9+8], 
           INIT[355*9+8], INIT[354*9+8], INIT[353*9+8], INIT[352*9+8], 
           INIT[351*9+8], INIT[350*9+8], INIT[349*9+8], INIT[348*9+8], 
           INIT[347*9+8], INIT[346*9+8], INIT[345*9+8], INIT[344*9+8], 
           INIT[343*9+8], INIT[342*9+8], INIT[341*9+8], INIT[340*9+8], 
           INIT[339*9+8], INIT[338*9+8], INIT[337*9+8], INIT[336*9+8], 
           INIT[335*9+8], INIT[334*9+8], INIT[333*9+8], INIT[332*9+8], 
           INIT[331*9+8], INIT[330*9+8], INIT[329*9+8], INIT[328*9+8], 
           INIT[327*9+8], INIT[326*9+8], INIT[325*9+8], INIT[324*9+8], 
           INIT[323*9+8], INIT[322*9+8], INIT[321*9+8], INIT[320*9+8], 
           INIT[319*9+8], INIT[318*9+8], INIT[317*9+8], INIT[316*9+8], 
           INIT[315*9+8], INIT[314*9+8], INIT[313*9+8], INIT[312*9+8], 
           INIT[311*9+8], INIT[310*9+8], INIT[309*9+8], INIT[308*9+8], 
           INIT[307*9+8], INIT[306*9+8], INIT[305*9+8], INIT[304*9+8], 
           INIT[303*9+8], INIT[302*9+8], INIT[301*9+8], INIT[300*9+8], 
           INIT[299*9+8], INIT[298*9+8], INIT[297*9+8], INIT[296*9+8], 
           INIT[295*9+8], INIT[294*9+8], INIT[293*9+8], INIT[292*9+8], 
           INIT[291*9+8], INIT[290*9+8], INIT[289*9+8], INIT[288*9+8], 
           INIT[287*9+8], INIT[286*9+8], INIT[285*9+8], INIT[284*9+8], 
           INIT[283*9+8], INIT[282*9+8], INIT[281*9+8], INIT[280*9+8], 
           INIT[279*9+8], INIT[278*9+8], INIT[277*9+8], INIT[276*9+8], 
           INIT[275*9+8], INIT[274*9+8], INIT[273*9+8], INIT[272*9+8], 
           INIT[271*9+8], INIT[270*9+8], INIT[269*9+8], INIT[268*9+8], 
           INIT[267*9+8], INIT[266*9+8], INIT[265*9+8], INIT[264*9+8], 
           INIT[263*9+8], INIT[262*9+8], INIT[261*9+8], INIT[260*9+8], 
           INIT[259*9+8], INIT[258*9+8], INIT[257*9+8], INIT[256*9+8]}),
.INITP_02({INIT[767*9+8], INIT[766*9+8], INIT[765*9+8], INIT[764*9+8], 
           INIT[763*9+8], INIT[762*9+8], INIT[761*9+8], INIT[760*9+8], 
           INIT[759*9+8], INIT[758*9+8], INIT[757*9+8], INIT[756*9+8], 
           INIT[755*9+8], INIT[754*9+8], INIT[753*9+8], INIT[752*9+8], 
           INIT[751*9+8], INIT[750*9+8], INIT[749*9+8], INIT[748*9+8], 
           INIT[747*9+8], INIT[746*9+8], INIT[745*9+8], INIT[744*9+8], 
           INIT[743*9+8], INIT[742*9+8], INIT[741*9+8], INIT[740*9+8], 
           INIT[739*9+8], INIT[738*9+8], INIT[737*9+8], INIT[736*9+8], 
           INIT[735*9+8], INIT[734*9+8], INIT[733*9+8], INIT[732*9+8], 
           INIT[731*9+8], INIT[730*9+8], INIT[729*9+8], INIT[728*9+8], 
           INIT[727*9+8], INIT[726*9+8], INIT[725*9+8], INIT[724*9+8], 
           INIT[723*9+8], INIT[722*9+8], INIT[721*9+8], INIT[720*9+8], 
           INIT[719*9+8], INIT[718*9+8], INIT[717*9+8], INIT[716*9+8], 
           INIT[715*9+8], INIT[714*9+8], INIT[713*9+8], INIT[712*9+8], 
           INIT[711*9+8], INIT[710*9+8], INIT[709*9+8], INIT[708*9+8], 
           INIT[707*9+8], INIT[706*9+8], INIT[705*9+8], INIT[704*9+8], 
           INIT[703*9+8], INIT[702*9+8], INIT[701*9+8], INIT[700*9+8], 
           INIT[699*9+8], INIT[698*9+8], INIT[697*9+8], INIT[696*9+8], 
           INIT[695*9+8], INIT[694*9+8], INIT[693*9+8], INIT[692*9+8], 
           INIT[691*9+8], INIT[690*9+8], INIT[689*9+8], INIT[688*9+8], 
           INIT[687*9+8], INIT[686*9+8], INIT[685*9+8], INIT[684*9+8], 
           INIT[683*9+8], INIT[682*9+8], INIT[681*9+8], INIT[680*9+8], 
           INIT[679*9+8], INIT[678*9+8], INIT[677*9+8], INIT[676*9+8], 
           INIT[675*9+8], INIT[674*9+8], INIT[673*9+8], INIT[672*9+8], 
           INIT[671*9+8], INIT[670*9+8], INIT[669*9+8], INIT[668*9+8], 
           INIT[667*9+8], INIT[666*9+8], INIT[665*9+8], INIT[664*9+8], 
           INIT[663*9+8], INIT[662*9+8], INIT[661*9+8], INIT[660*9+8], 
           INIT[659*9+8], INIT[658*9+8], INIT[657*9+8], INIT[656*9+8], 
           INIT[655*9+8], INIT[654*9+8], INIT[653*9+8], INIT[652*9+8], 
           INIT[651*9+8], INIT[650*9+8], INIT[649*9+8], INIT[648*9+8], 
           INIT[647*9+8], INIT[646*9+8], INIT[645*9+8], INIT[644*9+8], 
           INIT[643*9+8], INIT[642*9+8], INIT[641*9+8], INIT[640*9+8], 
           INIT[639*9+8], INIT[638*9+8], INIT[637*9+8], INIT[636*9+8], 
           INIT[635*9+8], INIT[634*9+8], INIT[633*9+8], INIT[632*9+8], 
           INIT[631*9+8], INIT[630*9+8], INIT[629*9+8], INIT[628*9+8], 
           INIT[627*9+8], INIT[626*9+8], INIT[625*9+8], INIT[624*9+8], 
           INIT[623*9+8], INIT[622*9+8], INIT[621*9+8], INIT[620*9+8], 
           INIT[619*9+8], INIT[618*9+8], INIT[617*9+8], INIT[616*9+8], 
           INIT[615*9+8], INIT[614*9+8], INIT[613*9+8], INIT[612*9+8], 
           INIT[611*9+8], INIT[610*9+8], INIT[609*9+8], INIT[608*9+8], 
           INIT[607*9+8], INIT[606*9+8], INIT[605*9+8], INIT[604*9+8], 
           INIT[603*9+8], INIT[602*9+8], INIT[601*9+8], INIT[600*9+8], 
           INIT[599*9+8], INIT[598*9+8], INIT[597*9+8], INIT[596*9+8], 
           INIT[595*9+8], INIT[594*9+8], INIT[593*9+8], INIT[592*9+8], 
           INIT[591*9+8], INIT[590*9+8], INIT[589*9+8], INIT[588*9+8], 
           INIT[587*9+8], INIT[586*9+8], INIT[585*9+8], INIT[584*9+8], 
           INIT[583*9+8], INIT[582*9+8], INIT[581*9+8], INIT[580*9+8], 
           INIT[579*9+8], INIT[578*9+8], INIT[577*9+8], INIT[576*9+8], 
           INIT[575*9+8], INIT[574*9+8], INIT[573*9+8], INIT[572*9+8], 
           INIT[571*9+8], INIT[570*9+8], INIT[569*9+8], INIT[568*9+8], 
           INIT[567*9+8], INIT[566*9+8], INIT[565*9+8], INIT[564*9+8], 
           INIT[563*9+8], INIT[562*9+8], INIT[561*9+8], INIT[560*9+8], 
           INIT[559*9+8], INIT[558*9+8], INIT[557*9+8], INIT[556*9+8], 
           INIT[555*9+8], INIT[554*9+8], INIT[553*9+8], INIT[552*9+8], 
           INIT[551*9+8], INIT[550*9+8], INIT[549*9+8], INIT[548*9+8], 
           INIT[547*9+8], INIT[546*9+8], INIT[545*9+8], INIT[544*9+8], 
           INIT[543*9+8], INIT[542*9+8], INIT[541*9+8], INIT[540*9+8], 
           INIT[539*9+8], INIT[538*9+8], INIT[537*9+8], INIT[536*9+8], 
           INIT[535*9+8], INIT[534*9+8], INIT[533*9+8], INIT[532*9+8], 
           INIT[531*9+8], INIT[530*9+8], INIT[529*9+8], INIT[528*9+8], 
           INIT[527*9+8], INIT[526*9+8], INIT[525*9+8], INIT[524*9+8], 
           INIT[523*9+8], INIT[522*9+8], INIT[521*9+8], INIT[520*9+8], 
           INIT[519*9+8], INIT[518*9+8], INIT[517*9+8], INIT[516*9+8], 
           INIT[515*9+8], INIT[514*9+8], INIT[513*9+8], INIT[512*9+8]}),
.INITP_03({INIT[1023*9+8], INIT[1022*9+8], INIT[1021*9+8], INIT[1020*9+8], 
           INIT[1019*9+8], INIT[1018*9+8], INIT[1017*9+8], INIT[1016*9+8], 
           INIT[1015*9+8], INIT[1014*9+8], INIT[1013*9+8], INIT[1012*9+8], 
           INIT[1011*9+8], INIT[1010*9+8], INIT[1009*9+8], INIT[1008*9+8], 
           INIT[1007*9+8], INIT[1006*9+8], INIT[1005*9+8], INIT[1004*9+8], 
           INIT[1003*9+8], INIT[1002*9+8], INIT[1001*9+8], INIT[1000*9+8], 
           INIT[999*9+8], INIT[998*9+8], INIT[997*9+8], INIT[996*9+8], 
           INIT[995*9+8], INIT[994*9+8], INIT[993*9+8], INIT[992*9+8], 
           INIT[991*9+8], INIT[990*9+8], INIT[989*9+8], INIT[988*9+8], 
           INIT[987*9+8], INIT[986*9+8], INIT[985*9+8], INIT[984*9+8], 
           INIT[983*9+8], INIT[982*9+8], INIT[981*9+8], INIT[980*9+8], 
           INIT[979*9+8], INIT[978*9+8], INIT[977*9+8], INIT[976*9+8], 
           INIT[975*9+8], INIT[974*9+8], INIT[973*9+8], INIT[972*9+8], 
           INIT[971*9+8], INIT[970*9+8], INIT[969*9+8], INIT[968*9+8], 
           INIT[967*9+8], INIT[966*9+8], INIT[965*9+8], INIT[964*9+8], 
           INIT[963*9+8], INIT[962*9+8], INIT[961*9+8], INIT[960*9+8], 
           INIT[959*9+8], INIT[958*9+8], INIT[957*9+8], INIT[956*9+8], 
           INIT[955*9+8], INIT[954*9+8], INIT[953*9+8], INIT[952*9+8], 
           INIT[951*9+8], INIT[950*9+8], INIT[949*9+8], INIT[948*9+8], 
           INIT[947*9+8], INIT[946*9+8], INIT[945*9+8], INIT[944*9+8], 
           INIT[943*9+8], INIT[942*9+8], INIT[941*9+8], INIT[940*9+8], 
           INIT[939*9+8], INIT[938*9+8], INIT[937*9+8], INIT[936*9+8], 
           INIT[935*9+8], INIT[934*9+8], INIT[933*9+8], INIT[932*9+8], 
           INIT[931*9+8], INIT[930*9+8], INIT[929*9+8], INIT[928*9+8], 
           INIT[927*9+8], INIT[926*9+8], INIT[925*9+8], INIT[924*9+8], 
           INIT[923*9+8], INIT[922*9+8], INIT[921*9+8], INIT[920*9+8], 
           INIT[919*9+8], INIT[918*9+8], INIT[917*9+8], INIT[916*9+8], 
           INIT[915*9+8], INIT[914*9+8], INIT[913*9+8], INIT[912*9+8], 
           INIT[911*9+8], INIT[910*9+8], INIT[909*9+8], INIT[908*9+8], 
           INIT[907*9+8], INIT[906*9+8], INIT[905*9+8], INIT[904*9+8], 
           INIT[903*9+8], INIT[902*9+8], INIT[901*9+8], INIT[900*9+8], 
           INIT[899*9+8], INIT[898*9+8], INIT[897*9+8], INIT[896*9+8], 
           INIT[895*9+8], INIT[894*9+8], INIT[893*9+8], INIT[892*9+8], 
           INIT[891*9+8], INIT[890*9+8], INIT[889*9+8], INIT[888*9+8], 
           INIT[887*9+8], INIT[886*9+8], INIT[885*9+8], INIT[884*9+8], 
           INIT[883*9+8], INIT[882*9+8], INIT[881*9+8], INIT[880*9+8], 
           INIT[879*9+8], INIT[878*9+8], INIT[877*9+8], INIT[876*9+8], 
           INIT[875*9+8], INIT[874*9+8], INIT[873*9+8], INIT[872*9+8], 
           INIT[871*9+8], INIT[870*9+8], INIT[869*9+8], INIT[868*9+8], 
           INIT[867*9+8], INIT[866*9+8], INIT[865*9+8], INIT[864*9+8], 
           INIT[863*9+8], INIT[862*9+8], INIT[861*9+8], INIT[860*9+8], 
           INIT[859*9+8], INIT[858*9+8], INIT[857*9+8], INIT[856*9+8], 
           INIT[855*9+8], INIT[854*9+8], INIT[853*9+8], INIT[852*9+8], 
           INIT[851*9+8], INIT[850*9+8], INIT[849*9+8], INIT[848*9+8], 
           INIT[847*9+8], INIT[846*9+8], INIT[845*9+8], INIT[844*9+8], 
           INIT[843*9+8], INIT[842*9+8], INIT[841*9+8], INIT[840*9+8], 
           INIT[839*9+8], INIT[838*9+8], INIT[837*9+8], INIT[836*9+8], 
           INIT[835*9+8], INIT[834*9+8], INIT[833*9+8], INIT[832*9+8], 
           INIT[831*9+8], INIT[830*9+8], INIT[829*9+8], INIT[828*9+8], 
           INIT[827*9+8], INIT[826*9+8], INIT[825*9+8], INIT[824*9+8], 
           INIT[823*9+8], INIT[822*9+8], INIT[821*9+8], INIT[820*9+8], 
           INIT[819*9+8], INIT[818*9+8], INIT[817*9+8], INIT[816*9+8], 
           INIT[815*9+8], INIT[814*9+8], INIT[813*9+8], INIT[812*9+8], 
           INIT[811*9+8], INIT[810*9+8], INIT[809*9+8], INIT[808*9+8], 
           INIT[807*9+8], INIT[806*9+8], INIT[805*9+8], INIT[804*9+8], 
           INIT[803*9+8], INIT[802*9+8], INIT[801*9+8], INIT[800*9+8], 
           INIT[799*9+8], INIT[798*9+8], INIT[797*9+8], INIT[796*9+8], 
           INIT[795*9+8], INIT[794*9+8], INIT[793*9+8], INIT[792*9+8], 
           INIT[791*9+8], INIT[790*9+8], INIT[789*9+8], INIT[788*9+8], 
           INIT[787*9+8], INIT[786*9+8], INIT[785*9+8], INIT[784*9+8], 
           INIT[783*9+8], INIT[782*9+8], INIT[781*9+8], INIT[780*9+8], 
           INIT[779*9+8], INIT[778*9+8], INIT[777*9+8], INIT[776*9+8], 
           INIT[775*9+8], INIT[774*9+8], INIT[773*9+8], INIT[772*9+8], 
           INIT[771*9+8], INIT[770*9+8], INIT[769*9+8], INIT[768*9+8]}),
.INITP_04({INIT[1279*9+8], INIT[1278*9+8], INIT[1277*9+8], INIT[1276*9+8], 
           INIT[1275*9+8], INIT[1274*9+8], INIT[1273*9+8], INIT[1272*9+8], 
           INIT[1271*9+8], INIT[1270*9+8], INIT[1269*9+8], INIT[1268*9+8], 
           INIT[1267*9+8], INIT[1266*9+8], INIT[1265*9+8], INIT[1264*9+8], 
           INIT[1263*9+8], INIT[1262*9+8], INIT[1261*9+8], INIT[1260*9+8], 
           INIT[1259*9+8], INIT[1258*9+8], INIT[1257*9+8], INIT[1256*9+8], 
           INIT[1255*9+8], INIT[1254*9+8], INIT[1253*9+8], INIT[1252*9+8], 
           INIT[1251*9+8], INIT[1250*9+8], INIT[1249*9+8], INIT[1248*9+8], 
           INIT[1247*9+8], INIT[1246*9+8], INIT[1245*9+8], INIT[1244*9+8], 
           INIT[1243*9+8], INIT[1242*9+8], INIT[1241*9+8], INIT[1240*9+8], 
           INIT[1239*9+8], INIT[1238*9+8], INIT[1237*9+8], INIT[1236*9+8], 
           INIT[1235*9+8], INIT[1234*9+8], INIT[1233*9+8], INIT[1232*9+8], 
           INIT[1231*9+8], INIT[1230*9+8], INIT[1229*9+8], INIT[1228*9+8], 
           INIT[1227*9+8], INIT[1226*9+8], INIT[1225*9+8], INIT[1224*9+8], 
           INIT[1223*9+8], INIT[1222*9+8], INIT[1221*9+8], INIT[1220*9+8], 
           INIT[1219*9+8], INIT[1218*9+8], INIT[1217*9+8], INIT[1216*9+8], 
           INIT[1215*9+8], INIT[1214*9+8], INIT[1213*9+8], INIT[1212*9+8], 
           INIT[1211*9+8], INIT[1210*9+8], INIT[1209*9+8], INIT[1208*9+8], 
           INIT[1207*9+8], INIT[1206*9+8], INIT[1205*9+8], INIT[1204*9+8], 
           INIT[1203*9+8], INIT[1202*9+8], INIT[1201*9+8], INIT[1200*9+8], 
           INIT[1199*9+8], INIT[1198*9+8], INIT[1197*9+8], INIT[1196*9+8], 
           INIT[1195*9+8], INIT[1194*9+8], INIT[1193*9+8], INIT[1192*9+8], 
           INIT[1191*9+8], INIT[1190*9+8], INIT[1189*9+8], INIT[1188*9+8], 
           INIT[1187*9+8], INIT[1186*9+8], INIT[1185*9+8], INIT[1184*9+8], 
           INIT[1183*9+8], INIT[1182*9+8], INIT[1181*9+8], INIT[1180*9+8], 
           INIT[1179*9+8], INIT[1178*9+8], INIT[1177*9+8], INIT[1176*9+8], 
           INIT[1175*9+8], INIT[1174*9+8], INIT[1173*9+8], INIT[1172*9+8], 
           INIT[1171*9+8], INIT[1170*9+8], INIT[1169*9+8], INIT[1168*9+8], 
           INIT[1167*9+8], INIT[1166*9+8], INIT[1165*9+8], INIT[1164*9+8], 
           INIT[1163*9+8], INIT[1162*9+8], INIT[1161*9+8], INIT[1160*9+8], 
           INIT[1159*9+8], INIT[1158*9+8], INIT[1157*9+8], INIT[1156*9+8], 
           INIT[1155*9+8], INIT[1154*9+8], INIT[1153*9+8], INIT[1152*9+8], 
           INIT[1151*9+8], INIT[1150*9+8], INIT[1149*9+8], INIT[1148*9+8], 
           INIT[1147*9+8], INIT[1146*9+8], INIT[1145*9+8], INIT[1144*9+8], 
           INIT[1143*9+8], INIT[1142*9+8], INIT[1141*9+8], INIT[1140*9+8], 
           INIT[1139*9+8], INIT[1138*9+8], INIT[1137*9+8], INIT[1136*9+8], 
           INIT[1135*9+8], INIT[1134*9+8], INIT[1133*9+8], INIT[1132*9+8], 
           INIT[1131*9+8], INIT[1130*9+8], INIT[1129*9+8], INIT[1128*9+8], 
           INIT[1127*9+8], INIT[1126*9+8], INIT[1125*9+8], INIT[1124*9+8], 
           INIT[1123*9+8], INIT[1122*9+8], INIT[1121*9+8], INIT[1120*9+8], 
           INIT[1119*9+8], INIT[1118*9+8], INIT[1117*9+8], INIT[1116*9+8], 
           INIT[1115*9+8], INIT[1114*9+8], INIT[1113*9+8], INIT[1112*9+8], 
           INIT[1111*9+8], INIT[1110*9+8], INIT[1109*9+8], INIT[1108*9+8], 
           INIT[1107*9+8], INIT[1106*9+8], INIT[1105*9+8], INIT[1104*9+8], 
           INIT[1103*9+8], INIT[1102*9+8], INIT[1101*9+8], INIT[1100*9+8], 
           INIT[1099*9+8], INIT[1098*9+8], INIT[1097*9+8], INIT[1096*9+8], 
           INIT[1095*9+8], INIT[1094*9+8], INIT[1093*9+8], INIT[1092*9+8], 
           INIT[1091*9+8], INIT[1090*9+8], INIT[1089*9+8], INIT[1088*9+8], 
           INIT[1087*9+8], INIT[1086*9+8], INIT[1085*9+8], INIT[1084*9+8], 
           INIT[1083*9+8], INIT[1082*9+8], INIT[1081*9+8], INIT[1080*9+8], 
           INIT[1079*9+8], INIT[1078*9+8], INIT[1077*9+8], INIT[1076*9+8], 
           INIT[1075*9+8], INIT[1074*9+8], INIT[1073*9+8], INIT[1072*9+8], 
           INIT[1071*9+8], INIT[1070*9+8], INIT[1069*9+8], INIT[1068*9+8], 
           INIT[1067*9+8], INIT[1066*9+8], INIT[1065*9+8], INIT[1064*9+8], 
           INIT[1063*9+8], INIT[1062*9+8], INIT[1061*9+8], INIT[1060*9+8], 
           INIT[1059*9+8], INIT[1058*9+8], INIT[1057*9+8], INIT[1056*9+8], 
           INIT[1055*9+8], INIT[1054*9+8], INIT[1053*9+8], INIT[1052*9+8], 
           INIT[1051*9+8], INIT[1050*9+8], INIT[1049*9+8], INIT[1048*9+8], 
           INIT[1047*9+8], INIT[1046*9+8], INIT[1045*9+8], INIT[1044*9+8], 
           INIT[1043*9+8], INIT[1042*9+8], INIT[1041*9+8], INIT[1040*9+8], 
           INIT[1039*9+8], INIT[1038*9+8], INIT[1037*9+8], INIT[1036*9+8], 
           INIT[1035*9+8], INIT[1034*9+8], INIT[1033*9+8], INIT[1032*9+8], 
           INIT[1031*9+8], INIT[1030*9+8], INIT[1029*9+8], INIT[1028*9+8], 
           INIT[1027*9+8], INIT[1026*9+8], INIT[1025*9+8], INIT[1024*9+8]}),
.INITP_05({INIT[1535*9+8], INIT[1534*9+8], INIT[1533*9+8], INIT[1532*9+8], 
           INIT[1531*9+8], INIT[1530*9+8], INIT[1529*9+8], INIT[1528*9+8], 
           INIT[1527*9+8], INIT[1526*9+8], INIT[1525*9+8], INIT[1524*9+8], 
           INIT[1523*9+8], INIT[1522*9+8], INIT[1521*9+8], INIT[1520*9+8], 
           INIT[1519*9+8], INIT[1518*9+8], INIT[1517*9+8], INIT[1516*9+8], 
           INIT[1515*9+8], INIT[1514*9+8], INIT[1513*9+8], INIT[1512*9+8], 
           INIT[1511*9+8], INIT[1510*9+8], INIT[1509*9+8], INIT[1508*9+8], 
           INIT[1507*9+8], INIT[1506*9+8], INIT[1505*9+8], INIT[1504*9+8], 
           INIT[1503*9+8], INIT[1502*9+8], INIT[1501*9+8], INIT[1500*9+8], 
           INIT[1499*9+8], INIT[1498*9+8], INIT[1497*9+8], INIT[1496*9+8], 
           INIT[1495*9+8], INIT[1494*9+8], INIT[1493*9+8], INIT[1492*9+8], 
           INIT[1491*9+8], INIT[1490*9+8], INIT[1489*9+8], INIT[1488*9+8], 
           INIT[1487*9+8], INIT[1486*9+8], INIT[1485*9+8], INIT[1484*9+8], 
           INIT[1483*9+8], INIT[1482*9+8], INIT[1481*9+8], INIT[1480*9+8], 
           INIT[1479*9+8], INIT[1478*9+8], INIT[1477*9+8], INIT[1476*9+8], 
           INIT[1475*9+8], INIT[1474*9+8], INIT[1473*9+8], INIT[1472*9+8], 
           INIT[1471*9+8], INIT[1470*9+8], INIT[1469*9+8], INIT[1468*9+8], 
           INIT[1467*9+8], INIT[1466*9+8], INIT[1465*9+8], INIT[1464*9+8], 
           INIT[1463*9+8], INIT[1462*9+8], INIT[1461*9+8], INIT[1460*9+8], 
           INIT[1459*9+8], INIT[1458*9+8], INIT[1457*9+8], INIT[1456*9+8], 
           INIT[1455*9+8], INIT[1454*9+8], INIT[1453*9+8], INIT[1452*9+8], 
           INIT[1451*9+8], INIT[1450*9+8], INIT[1449*9+8], INIT[1448*9+8], 
           INIT[1447*9+8], INIT[1446*9+8], INIT[1445*9+8], INIT[1444*9+8], 
           INIT[1443*9+8], INIT[1442*9+8], INIT[1441*9+8], INIT[1440*9+8], 
           INIT[1439*9+8], INIT[1438*9+8], INIT[1437*9+8], INIT[1436*9+8], 
           INIT[1435*9+8], INIT[1434*9+8], INIT[1433*9+8], INIT[1432*9+8], 
           INIT[1431*9+8], INIT[1430*9+8], INIT[1429*9+8], INIT[1428*9+8], 
           INIT[1427*9+8], INIT[1426*9+8], INIT[1425*9+8], INIT[1424*9+8], 
           INIT[1423*9+8], INIT[1422*9+8], INIT[1421*9+8], INIT[1420*9+8], 
           INIT[1419*9+8], INIT[1418*9+8], INIT[1417*9+8], INIT[1416*9+8], 
           INIT[1415*9+8], INIT[1414*9+8], INIT[1413*9+8], INIT[1412*9+8], 
           INIT[1411*9+8], INIT[1410*9+8], INIT[1409*9+8], INIT[1408*9+8], 
           INIT[1407*9+8], INIT[1406*9+8], INIT[1405*9+8], INIT[1404*9+8], 
           INIT[1403*9+8], INIT[1402*9+8], INIT[1401*9+8], INIT[1400*9+8], 
           INIT[1399*9+8], INIT[1398*9+8], INIT[1397*9+8], INIT[1396*9+8], 
           INIT[1395*9+8], INIT[1394*9+8], INIT[1393*9+8], INIT[1392*9+8], 
           INIT[1391*9+8], INIT[1390*9+8], INIT[1389*9+8], INIT[1388*9+8], 
           INIT[1387*9+8], INIT[1386*9+8], INIT[1385*9+8], INIT[1384*9+8], 
           INIT[1383*9+8], INIT[1382*9+8], INIT[1381*9+8], INIT[1380*9+8], 
           INIT[1379*9+8], INIT[1378*9+8], INIT[1377*9+8], INIT[1376*9+8], 
           INIT[1375*9+8], INIT[1374*9+8], INIT[1373*9+8], INIT[1372*9+8], 
           INIT[1371*9+8], INIT[1370*9+8], INIT[1369*9+8], INIT[1368*9+8], 
           INIT[1367*9+8], INIT[1366*9+8], INIT[1365*9+8], INIT[1364*9+8], 
           INIT[1363*9+8], INIT[1362*9+8], INIT[1361*9+8], INIT[1360*9+8], 
           INIT[1359*9+8], INIT[1358*9+8], INIT[1357*9+8], INIT[1356*9+8], 
           INIT[1355*9+8], INIT[1354*9+8], INIT[1353*9+8], INIT[1352*9+8], 
           INIT[1351*9+8], INIT[1350*9+8], INIT[1349*9+8], INIT[1348*9+8], 
           INIT[1347*9+8], INIT[1346*9+8], INIT[1345*9+8], INIT[1344*9+8], 
           INIT[1343*9+8], INIT[1342*9+8], INIT[1341*9+8], INIT[1340*9+8], 
           INIT[1339*9+8], INIT[1338*9+8], INIT[1337*9+8], INIT[1336*9+8], 
           INIT[1335*9+8], INIT[1334*9+8], INIT[1333*9+8], INIT[1332*9+8], 
           INIT[1331*9+8], INIT[1330*9+8], INIT[1329*9+8], INIT[1328*9+8], 
           INIT[1327*9+8], INIT[1326*9+8], INIT[1325*9+8], INIT[1324*9+8], 
           INIT[1323*9+8], INIT[1322*9+8], INIT[1321*9+8], INIT[1320*9+8], 
           INIT[1319*9+8], INIT[1318*9+8], INIT[1317*9+8], INIT[1316*9+8], 
           INIT[1315*9+8], INIT[1314*9+8], INIT[1313*9+8], INIT[1312*9+8], 
           INIT[1311*9+8], INIT[1310*9+8], INIT[1309*9+8], INIT[1308*9+8], 
           INIT[1307*9+8], INIT[1306*9+8], INIT[1305*9+8], INIT[1304*9+8], 
           INIT[1303*9+8], INIT[1302*9+8], INIT[1301*9+8], INIT[1300*9+8], 
           INIT[1299*9+8], INIT[1298*9+8], INIT[1297*9+8], INIT[1296*9+8], 
           INIT[1295*9+8], INIT[1294*9+8], INIT[1293*9+8], INIT[1292*9+8], 
           INIT[1291*9+8], INIT[1290*9+8], INIT[1289*9+8], INIT[1288*9+8], 
           INIT[1287*9+8], INIT[1286*9+8], INIT[1285*9+8], INIT[1284*9+8], 
           INIT[1283*9+8], INIT[1282*9+8], INIT[1281*9+8], INIT[1280*9+8]}),
.INITP_06({INIT[1791*9+8], INIT[1790*9+8], INIT[1789*9+8], INIT[1788*9+8], 
           INIT[1787*9+8], INIT[1786*9+8], INIT[1785*9+8], INIT[1784*9+8], 
           INIT[1783*9+8], INIT[1782*9+8], INIT[1781*9+8], INIT[1780*9+8], 
           INIT[1779*9+8], INIT[1778*9+8], INIT[1777*9+8], INIT[1776*9+8], 
           INIT[1775*9+8], INIT[1774*9+8], INIT[1773*9+8], INIT[1772*9+8], 
           INIT[1771*9+8], INIT[1770*9+8], INIT[1769*9+8], INIT[1768*9+8], 
           INIT[1767*9+8], INIT[1766*9+8], INIT[1765*9+8], INIT[1764*9+8], 
           INIT[1763*9+8], INIT[1762*9+8], INIT[1761*9+8], INIT[1760*9+8], 
           INIT[1759*9+8], INIT[1758*9+8], INIT[1757*9+8], INIT[1756*9+8], 
           INIT[1755*9+8], INIT[1754*9+8], INIT[1753*9+8], INIT[1752*9+8], 
           INIT[1751*9+8], INIT[1750*9+8], INIT[1749*9+8], INIT[1748*9+8], 
           INIT[1747*9+8], INIT[1746*9+8], INIT[1745*9+8], INIT[1744*9+8], 
           INIT[1743*9+8], INIT[1742*9+8], INIT[1741*9+8], INIT[1740*9+8], 
           INIT[1739*9+8], INIT[1738*9+8], INIT[1737*9+8], INIT[1736*9+8], 
           INIT[1735*9+8], INIT[1734*9+8], INIT[1733*9+8], INIT[1732*9+8], 
           INIT[1731*9+8], INIT[1730*9+8], INIT[1729*9+8], INIT[1728*9+8], 
           INIT[1727*9+8], INIT[1726*9+8], INIT[1725*9+8], INIT[1724*9+8], 
           INIT[1723*9+8], INIT[1722*9+8], INIT[1721*9+8], INIT[1720*9+8], 
           INIT[1719*9+8], INIT[1718*9+8], INIT[1717*9+8], INIT[1716*9+8], 
           INIT[1715*9+8], INIT[1714*9+8], INIT[1713*9+8], INIT[1712*9+8], 
           INIT[1711*9+8], INIT[1710*9+8], INIT[1709*9+8], INIT[1708*9+8], 
           INIT[1707*9+8], INIT[1706*9+8], INIT[1705*9+8], INIT[1704*9+8], 
           INIT[1703*9+8], INIT[1702*9+8], INIT[1701*9+8], INIT[1700*9+8], 
           INIT[1699*9+8], INIT[1698*9+8], INIT[1697*9+8], INIT[1696*9+8], 
           INIT[1695*9+8], INIT[1694*9+8], INIT[1693*9+8], INIT[1692*9+8], 
           INIT[1691*9+8], INIT[1690*9+8], INIT[1689*9+8], INIT[1688*9+8], 
           INIT[1687*9+8], INIT[1686*9+8], INIT[1685*9+8], INIT[1684*9+8], 
           INIT[1683*9+8], INIT[1682*9+8], INIT[1681*9+8], INIT[1680*9+8], 
           INIT[1679*9+8], INIT[1678*9+8], INIT[1677*9+8], INIT[1676*9+8], 
           INIT[1675*9+8], INIT[1674*9+8], INIT[1673*9+8], INIT[1672*9+8], 
           INIT[1671*9+8], INIT[1670*9+8], INIT[1669*9+8], INIT[1668*9+8], 
           INIT[1667*9+8], INIT[1666*9+8], INIT[1665*9+8], INIT[1664*9+8], 
           INIT[1663*9+8], INIT[1662*9+8], INIT[1661*9+8], INIT[1660*9+8], 
           INIT[1659*9+8], INIT[1658*9+8], INIT[1657*9+8], INIT[1656*9+8], 
           INIT[1655*9+8], INIT[1654*9+8], INIT[1653*9+8], INIT[1652*9+8], 
           INIT[1651*9+8], INIT[1650*9+8], INIT[1649*9+8], INIT[1648*9+8], 
           INIT[1647*9+8], INIT[1646*9+8], INIT[1645*9+8], INIT[1644*9+8], 
           INIT[1643*9+8], INIT[1642*9+8], INIT[1641*9+8], INIT[1640*9+8], 
           INIT[1639*9+8], INIT[1638*9+8], INIT[1637*9+8], INIT[1636*9+8], 
           INIT[1635*9+8], INIT[1634*9+8], INIT[1633*9+8], INIT[1632*9+8], 
           INIT[1631*9+8], INIT[1630*9+8], INIT[1629*9+8], INIT[1628*9+8], 
           INIT[1627*9+8], INIT[1626*9+8], INIT[1625*9+8], INIT[1624*9+8], 
           INIT[1623*9+8], INIT[1622*9+8], INIT[1621*9+8], INIT[1620*9+8], 
           INIT[1619*9+8], INIT[1618*9+8], INIT[1617*9+8], INIT[1616*9+8], 
           INIT[1615*9+8], INIT[1614*9+8], INIT[1613*9+8], INIT[1612*9+8], 
           INIT[1611*9+8], INIT[1610*9+8], INIT[1609*9+8], INIT[1608*9+8], 
           INIT[1607*9+8], INIT[1606*9+8], INIT[1605*9+8], INIT[1604*9+8], 
           INIT[1603*9+8], INIT[1602*9+8], INIT[1601*9+8], INIT[1600*9+8], 
           INIT[1599*9+8], INIT[1598*9+8], INIT[1597*9+8], INIT[1596*9+8], 
           INIT[1595*9+8], INIT[1594*9+8], INIT[1593*9+8], INIT[1592*9+8], 
           INIT[1591*9+8], INIT[1590*9+8], INIT[1589*9+8], INIT[1588*9+8], 
           INIT[1587*9+8], INIT[1586*9+8], INIT[1585*9+8], INIT[1584*9+8], 
           INIT[1583*9+8], INIT[1582*9+8], INIT[1581*9+8], INIT[1580*9+8], 
           INIT[1579*9+8], INIT[1578*9+8], INIT[1577*9+8], INIT[1576*9+8], 
           INIT[1575*9+8], INIT[1574*9+8], INIT[1573*9+8], INIT[1572*9+8], 
           INIT[1571*9+8], INIT[1570*9+8], INIT[1569*9+8], INIT[1568*9+8], 
           INIT[1567*9+8], INIT[1566*9+8], INIT[1565*9+8], INIT[1564*9+8], 
           INIT[1563*9+8], INIT[1562*9+8], INIT[1561*9+8], INIT[1560*9+8], 
           INIT[1559*9+8], INIT[1558*9+8], INIT[1557*9+8], INIT[1556*9+8], 
           INIT[1555*9+8], INIT[1554*9+8], INIT[1553*9+8], INIT[1552*9+8], 
           INIT[1551*9+8], INIT[1550*9+8], INIT[1549*9+8], INIT[1548*9+8], 
           INIT[1547*9+8], INIT[1546*9+8], INIT[1545*9+8], INIT[1544*9+8], 
           INIT[1543*9+8], INIT[1542*9+8], INIT[1541*9+8], INIT[1540*9+8], 
           INIT[1539*9+8], INIT[1538*9+8], INIT[1537*9+8], INIT[1536*9+8]}),
.INITP_07({INIT[2047*9+8], INIT[2046*9+8], INIT[2045*9+8], INIT[2044*9+8], 
           INIT[2043*9+8], INIT[2042*9+8], INIT[2041*9+8], INIT[2040*9+8], 
           INIT[2039*9+8], INIT[2038*9+8], INIT[2037*9+8], INIT[2036*9+8], 
           INIT[2035*9+8], INIT[2034*9+8], INIT[2033*9+8], INIT[2032*9+8], 
           INIT[2031*9+8], INIT[2030*9+8], INIT[2029*9+8], INIT[2028*9+8], 
           INIT[2027*9+8], INIT[2026*9+8], INIT[2025*9+8], INIT[2024*9+8], 
           INIT[2023*9+8], INIT[2022*9+8], INIT[2021*9+8], INIT[2020*9+8], 
           INIT[2019*9+8], INIT[2018*9+8], INIT[2017*9+8], INIT[2016*9+8], 
           INIT[2015*9+8], INIT[2014*9+8], INIT[2013*9+8], INIT[2012*9+8], 
           INIT[2011*9+8], INIT[2010*9+8], INIT[2009*9+8], INIT[2008*9+8], 
           INIT[2007*9+8], INIT[2006*9+8], INIT[2005*9+8], INIT[2004*9+8], 
           INIT[2003*9+8], INIT[2002*9+8], INIT[2001*9+8], INIT[2000*9+8], 
           INIT[1999*9+8], INIT[1998*9+8], INIT[1997*9+8], INIT[1996*9+8], 
           INIT[1995*9+8], INIT[1994*9+8], INIT[1993*9+8], INIT[1992*9+8], 
           INIT[1991*9+8], INIT[1990*9+8], INIT[1989*9+8], INIT[1988*9+8], 
           INIT[1987*9+8], INIT[1986*9+8], INIT[1985*9+8], INIT[1984*9+8], 
           INIT[1983*9+8], INIT[1982*9+8], INIT[1981*9+8], INIT[1980*9+8], 
           INIT[1979*9+8], INIT[1978*9+8], INIT[1977*9+8], INIT[1976*9+8], 
           INIT[1975*9+8], INIT[1974*9+8], INIT[1973*9+8], INIT[1972*9+8], 
           INIT[1971*9+8], INIT[1970*9+8], INIT[1969*9+8], INIT[1968*9+8], 
           INIT[1967*9+8], INIT[1966*9+8], INIT[1965*9+8], INIT[1964*9+8], 
           INIT[1963*9+8], INIT[1962*9+8], INIT[1961*9+8], INIT[1960*9+8], 
           INIT[1959*9+8], INIT[1958*9+8], INIT[1957*9+8], INIT[1956*9+8], 
           INIT[1955*9+8], INIT[1954*9+8], INIT[1953*9+8], INIT[1952*9+8], 
           INIT[1951*9+8], INIT[1950*9+8], INIT[1949*9+8], INIT[1948*9+8], 
           INIT[1947*9+8], INIT[1946*9+8], INIT[1945*9+8], INIT[1944*9+8], 
           INIT[1943*9+8], INIT[1942*9+8], INIT[1941*9+8], INIT[1940*9+8], 
           INIT[1939*9+8], INIT[1938*9+8], INIT[1937*9+8], INIT[1936*9+8], 
           INIT[1935*9+8], INIT[1934*9+8], INIT[1933*9+8], INIT[1932*9+8], 
           INIT[1931*9+8], INIT[1930*9+8], INIT[1929*9+8], INIT[1928*9+8], 
           INIT[1927*9+8], INIT[1926*9+8], INIT[1925*9+8], INIT[1924*9+8], 
           INIT[1923*9+8], INIT[1922*9+8], INIT[1921*9+8], INIT[1920*9+8], 
           INIT[1919*9+8], INIT[1918*9+8], INIT[1917*9+8], INIT[1916*9+8], 
           INIT[1915*9+8], INIT[1914*9+8], INIT[1913*9+8], INIT[1912*9+8], 
           INIT[1911*9+8], INIT[1910*9+8], INIT[1909*9+8], INIT[1908*9+8], 
           INIT[1907*9+8], INIT[1906*9+8], INIT[1905*9+8], INIT[1904*9+8], 
           INIT[1903*9+8], INIT[1902*9+8], INIT[1901*9+8], INIT[1900*9+8], 
           INIT[1899*9+8], INIT[1898*9+8], INIT[1897*9+8], INIT[1896*9+8], 
           INIT[1895*9+8], INIT[1894*9+8], INIT[1893*9+8], INIT[1892*9+8], 
           INIT[1891*9+8], INIT[1890*9+8], INIT[1889*9+8], INIT[1888*9+8], 
           INIT[1887*9+8], INIT[1886*9+8], INIT[1885*9+8], INIT[1884*9+8], 
           INIT[1883*9+8], INIT[1882*9+8], INIT[1881*9+8], INIT[1880*9+8], 
           INIT[1879*9+8], INIT[1878*9+8], INIT[1877*9+8], INIT[1876*9+8], 
           INIT[1875*9+8], INIT[1874*9+8], INIT[1873*9+8], INIT[1872*9+8], 
           INIT[1871*9+8], INIT[1870*9+8], INIT[1869*9+8], INIT[1868*9+8], 
           INIT[1867*9+8], INIT[1866*9+8], INIT[1865*9+8], INIT[1864*9+8], 
           INIT[1863*9+8], INIT[1862*9+8], INIT[1861*9+8], INIT[1860*9+8], 
           INIT[1859*9+8], INIT[1858*9+8], INIT[1857*9+8], INIT[1856*9+8], 
           INIT[1855*9+8], INIT[1854*9+8], INIT[1853*9+8], INIT[1852*9+8], 
           INIT[1851*9+8], INIT[1850*9+8], INIT[1849*9+8], INIT[1848*9+8], 
           INIT[1847*9+8], INIT[1846*9+8], INIT[1845*9+8], INIT[1844*9+8], 
           INIT[1843*9+8], INIT[1842*9+8], INIT[1841*9+8], INIT[1840*9+8], 
           INIT[1839*9+8], INIT[1838*9+8], INIT[1837*9+8], INIT[1836*9+8], 
           INIT[1835*9+8], INIT[1834*9+8], INIT[1833*9+8], INIT[1832*9+8], 
           INIT[1831*9+8], INIT[1830*9+8], INIT[1829*9+8], INIT[1828*9+8], 
           INIT[1827*9+8], INIT[1826*9+8], INIT[1825*9+8], INIT[1824*9+8], 
           INIT[1823*9+8], INIT[1822*9+8], INIT[1821*9+8], INIT[1820*9+8], 
           INIT[1819*9+8], INIT[1818*9+8], INIT[1817*9+8], INIT[1816*9+8], 
           INIT[1815*9+8], INIT[1814*9+8], INIT[1813*9+8], INIT[1812*9+8], 
           INIT[1811*9+8], INIT[1810*9+8], INIT[1809*9+8], INIT[1808*9+8], 
           INIT[1807*9+8], INIT[1806*9+8], INIT[1805*9+8], INIT[1804*9+8], 
           INIT[1803*9+8], INIT[1802*9+8], INIT[1801*9+8], INIT[1800*9+8], 
           INIT[1799*9+8], INIT[1798*9+8], INIT[1797*9+8], INIT[1796*9+8], 
           INIT[1795*9+8], INIT[1794*9+8], INIT[1793*9+8], INIT[1792*9+8]}),
.INITP_08({INIT[2303*9+8], INIT[2302*9+8], INIT[2301*9+8], INIT[2300*9+8], 
           INIT[2299*9+8], INIT[2298*9+8], INIT[2297*9+8], INIT[2296*9+8], 
           INIT[2295*9+8], INIT[2294*9+8], INIT[2293*9+8], INIT[2292*9+8], 
           INIT[2291*9+8], INIT[2290*9+8], INIT[2289*9+8], INIT[2288*9+8], 
           INIT[2287*9+8], INIT[2286*9+8], INIT[2285*9+8], INIT[2284*9+8], 
           INIT[2283*9+8], INIT[2282*9+8], INIT[2281*9+8], INIT[2280*9+8], 
           INIT[2279*9+8], INIT[2278*9+8], INIT[2277*9+8], INIT[2276*9+8], 
           INIT[2275*9+8], INIT[2274*9+8], INIT[2273*9+8], INIT[2272*9+8], 
           INIT[2271*9+8], INIT[2270*9+8], INIT[2269*9+8], INIT[2268*9+8], 
           INIT[2267*9+8], INIT[2266*9+8], INIT[2265*9+8], INIT[2264*9+8], 
           INIT[2263*9+8], INIT[2262*9+8], INIT[2261*9+8], INIT[2260*9+8], 
           INIT[2259*9+8], INIT[2258*9+8], INIT[2257*9+8], INIT[2256*9+8], 
           INIT[2255*9+8], INIT[2254*9+8], INIT[2253*9+8], INIT[2252*9+8], 
           INIT[2251*9+8], INIT[2250*9+8], INIT[2249*9+8], INIT[2248*9+8], 
           INIT[2247*9+8], INIT[2246*9+8], INIT[2245*9+8], INIT[2244*9+8], 
           INIT[2243*9+8], INIT[2242*9+8], INIT[2241*9+8], INIT[2240*9+8], 
           INIT[2239*9+8], INIT[2238*9+8], INIT[2237*9+8], INIT[2236*9+8], 
           INIT[2235*9+8], INIT[2234*9+8], INIT[2233*9+8], INIT[2232*9+8], 
           INIT[2231*9+8], INIT[2230*9+8], INIT[2229*9+8], INIT[2228*9+8], 
           INIT[2227*9+8], INIT[2226*9+8], INIT[2225*9+8], INIT[2224*9+8], 
           INIT[2223*9+8], INIT[2222*9+8], INIT[2221*9+8], INIT[2220*9+8], 
           INIT[2219*9+8], INIT[2218*9+8], INIT[2217*9+8], INIT[2216*9+8], 
           INIT[2215*9+8], INIT[2214*9+8], INIT[2213*9+8], INIT[2212*9+8], 
           INIT[2211*9+8], INIT[2210*9+8], INIT[2209*9+8], INIT[2208*9+8], 
           INIT[2207*9+8], INIT[2206*9+8], INIT[2205*9+8], INIT[2204*9+8], 
           INIT[2203*9+8], INIT[2202*9+8], INIT[2201*9+8], INIT[2200*9+8], 
           INIT[2199*9+8], INIT[2198*9+8], INIT[2197*9+8], INIT[2196*9+8], 
           INIT[2195*9+8], INIT[2194*9+8], INIT[2193*9+8], INIT[2192*9+8], 
           INIT[2191*9+8], INIT[2190*9+8], INIT[2189*9+8], INIT[2188*9+8], 
           INIT[2187*9+8], INIT[2186*9+8], INIT[2185*9+8], INIT[2184*9+8], 
           INIT[2183*9+8], INIT[2182*9+8], INIT[2181*9+8], INIT[2180*9+8], 
           INIT[2179*9+8], INIT[2178*9+8], INIT[2177*9+8], INIT[2176*9+8], 
           INIT[2175*9+8], INIT[2174*9+8], INIT[2173*9+8], INIT[2172*9+8], 
           INIT[2171*9+8], INIT[2170*9+8], INIT[2169*9+8], INIT[2168*9+8], 
           INIT[2167*9+8], INIT[2166*9+8], INIT[2165*9+8], INIT[2164*9+8], 
           INIT[2163*9+8], INIT[2162*9+8], INIT[2161*9+8], INIT[2160*9+8], 
           INIT[2159*9+8], INIT[2158*9+8], INIT[2157*9+8], INIT[2156*9+8], 
           INIT[2155*9+8], INIT[2154*9+8], INIT[2153*9+8], INIT[2152*9+8], 
           INIT[2151*9+8], INIT[2150*9+8], INIT[2149*9+8], INIT[2148*9+8], 
           INIT[2147*9+8], INIT[2146*9+8], INIT[2145*9+8], INIT[2144*9+8], 
           INIT[2143*9+8], INIT[2142*9+8], INIT[2141*9+8], INIT[2140*9+8], 
           INIT[2139*9+8], INIT[2138*9+8], INIT[2137*9+8], INIT[2136*9+8], 
           INIT[2135*9+8], INIT[2134*9+8], INIT[2133*9+8], INIT[2132*9+8], 
           INIT[2131*9+8], INIT[2130*9+8], INIT[2129*9+8], INIT[2128*9+8], 
           INIT[2127*9+8], INIT[2126*9+8], INIT[2125*9+8], INIT[2124*9+8], 
           INIT[2123*9+8], INIT[2122*9+8], INIT[2121*9+8], INIT[2120*9+8], 
           INIT[2119*9+8], INIT[2118*9+8], INIT[2117*9+8], INIT[2116*9+8], 
           INIT[2115*9+8], INIT[2114*9+8], INIT[2113*9+8], INIT[2112*9+8], 
           INIT[2111*9+8], INIT[2110*9+8], INIT[2109*9+8], INIT[2108*9+8], 
           INIT[2107*9+8], INIT[2106*9+8], INIT[2105*9+8], INIT[2104*9+8], 
           INIT[2103*9+8], INIT[2102*9+8], INIT[2101*9+8], INIT[2100*9+8], 
           INIT[2099*9+8], INIT[2098*9+8], INIT[2097*9+8], INIT[2096*9+8], 
           INIT[2095*9+8], INIT[2094*9+8], INIT[2093*9+8], INIT[2092*9+8], 
           INIT[2091*9+8], INIT[2090*9+8], INIT[2089*9+8], INIT[2088*9+8], 
           INIT[2087*9+8], INIT[2086*9+8], INIT[2085*9+8], INIT[2084*9+8], 
           INIT[2083*9+8], INIT[2082*9+8], INIT[2081*9+8], INIT[2080*9+8], 
           INIT[2079*9+8], INIT[2078*9+8], INIT[2077*9+8], INIT[2076*9+8], 
           INIT[2075*9+8], INIT[2074*9+8], INIT[2073*9+8], INIT[2072*9+8], 
           INIT[2071*9+8], INIT[2070*9+8], INIT[2069*9+8], INIT[2068*9+8], 
           INIT[2067*9+8], INIT[2066*9+8], INIT[2065*9+8], INIT[2064*9+8], 
           INIT[2063*9+8], INIT[2062*9+8], INIT[2061*9+8], INIT[2060*9+8], 
           INIT[2059*9+8], INIT[2058*9+8], INIT[2057*9+8], INIT[2056*9+8], 
           INIT[2055*9+8], INIT[2054*9+8], INIT[2053*9+8], INIT[2052*9+8], 
           INIT[2051*9+8], INIT[2050*9+8], INIT[2049*9+8], INIT[2048*9+8]}),
.INITP_09({INIT[2559*9+8], INIT[2558*9+8], INIT[2557*9+8], INIT[2556*9+8], 
           INIT[2555*9+8], INIT[2554*9+8], INIT[2553*9+8], INIT[2552*9+8], 
           INIT[2551*9+8], INIT[2550*9+8], INIT[2549*9+8], INIT[2548*9+8], 
           INIT[2547*9+8], INIT[2546*9+8], INIT[2545*9+8], INIT[2544*9+8], 
           INIT[2543*9+8], INIT[2542*9+8], INIT[2541*9+8], INIT[2540*9+8], 
           INIT[2539*9+8], INIT[2538*9+8], INIT[2537*9+8], INIT[2536*9+8], 
           INIT[2535*9+8], INIT[2534*9+8], INIT[2533*9+8], INIT[2532*9+8], 
           INIT[2531*9+8], INIT[2530*9+8], INIT[2529*9+8], INIT[2528*9+8], 
           INIT[2527*9+8], INIT[2526*9+8], INIT[2525*9+8], INIT[2524*9+8], 
           INIT[2523*9+8], INIT[2522*9+8], INIT[2521*9+8], INIT[2520*9+8], 
           INIT[2519*9+8], INIT[2518*9+8], INIT[2517*9+8], INIT[2516*9+8], 
           INIT[2515*9+8], INIT[2514*9+8], INIT[2513*9+8], INIT[2512*9+8], 
           INIT[2511*9+8], INIT[2510*9+8], INIT[2509*9+8], INIT[2508*9+8], 
           INIT[2507*9+8], INIT[2506*9+8], INIT[2505*9+8], INIT[2504*9+8], 
           INIT[2503*9+8], INIT[2502*9+8], INIT[2501*9+8], INIT[2500*9+8], 
           INIT[2499*9+8], INIT[2498*9+8], INIT[2497*9+8], INIT[2496*9+8], 
           INIT[2495*9+8], INIT[2494*9+8], INIT[2493*9+8], INIT[2492*9+8], 
           INIT[2491*9+8], INIT[2490*9+8], INIT[2489*9+8], INIT[2488*9+8], 
           INIT[2487*9+8], INIT[2486*9+8], INIT[2485*9+8], INIT[2484*9+8], 
           INIT[2483*9+8], INIT[2482*9+8], INIT[2481*9+8], INIT[2480*9+8], 
           INIT[2479*9+8], INIT[2478*9+8], INIT[2477*9+8], INIT[2476*9+8], 
           INIT[2475*9+8], INIT[2474*9+8], INIT[2473*9+8], INIT[2472*9+8], 
           INIT[2471*9+8], INIT[2470*9+8], INIT[2469*9+8], INIT[2468*9+8], 
           INIT[2467*9+8], INIT[2466*9+8], INIT[2465*9+8], INIT[2464*9+8], 
           INIT[2463*9+8], INIT[2462*9+8], INIT[2461*9+8], INIT[2460*9+8], 
           INIT[2459*9+8], INIT[2458*9+8], INIT[2457*9+8], INIT[2456*9+8], 
           INIT[2455*9+8], INIT[2454*9+8], INIT[2453*9+8], INIT[2452*9+8], 
           INIT[2451*9+8], INIT[2450*9+8], INIT[2449*9+8], INIT[2448*9+8], 
           INIT[2447*9+8], INIT[2446*9+8], INIT[2445*9+8], INIT[2444*9+8], 
           INIT[2443*9+8], INIT[2442*9+8], INIT[2441*9+8], INIT[2440*9+8], 
           INIT[2439*9+8], INIT[2438*9+8], INIT[2437*9+8], INIT[2436*9+8], 
           INIT[2435*9+8], INIT[2434*9+8], INIT[2433*9+8], INIT[2432*9+8], 
           INIT[2431*9+8], INIT[2430*9+8], INIT[2429*9+8], INIT[2428*9+8], 
           INIT[2427*9+8], INIT[2426*9+8], INIT[2425*9+8], INIT[2424*9+8], 
           INIT[2423*9+8], INIT[2422*9+8], INIT[2421*9+8], INIT[2420*9+8], 
           INIT[2419*9+8], INIT[2418*9+8], INIT[2417*9+8], INIT[2416*9+8], 
           INIT[2415*9+8], INIT[2414*9+8], INIT[2413*9+8], INIT[2412*9+8], 
           INIT[2411*9+8], INIT[2410*9+8], INIT[2409*9+8], INIT[2408*9+8], 
           INIT[2407*9+8], INIT[2406*9+8], INIT[2405*9+8], INIT[2404*9+8], 
           INIT[2403*9+8], INIT[2402*9+8], INIT[2401*9+8], INIT[2400*9+8], 
           INIT[2399*9+8], INIT[2398*9+8], INIT[2397*9+8], INIT[2396*9+8], 
           INIT[2395*9+8], INIT[2394*9+8], INIT[2393*9+8], INIT[2392*9+8], 
           INIT[2391*9+8], INIT[2390*9+8], INIT[2389*9+8], INIT[2388*9+8], 
           INIT[2387*9+8], INIT[2386*9+8], INIT[2385*9+8], INIT[2384*9+8], 
           INIT[2383*9+8], INIT[2382*9+8], INIT[2381*9+8], INIT[2380*9+8], 
           INIT[2379*9+8], INIT[2378*9+8], INIT[2377*9+8], INIT[2376*9+8], 
           INIT[2375*9+8], INIT[2374*9+8], INIT[2373*9+8], INIT[2372*9+8], 
           INIT[2371*9+8], INIT[2370*9+8], INIT[2369*9+8], INIT[2368*9+8], 
           INIT[2367*9+8], INIT[2366*9+8], INIT[2365*9+8], INIT[2364*9+8], 
           INIT[2363*9+8], INIT[2362*9+8], INIT[2361*9+8], INIT[2360*9+8], 
           INIT[2359*9+8], INIT[2358*9+8], INIT[2357*9+8], INIT[2356*9+8], 
           INIT[2355*9+8], INIT[2354*9+8], INIT[2353*9+8], INIT[2352*9+8], 
           INIT[2351*9+8], INIT[2350*9+8], INIT[2349*9+8], INIT[2348*9+8], 
           INIT[2347*9+8], INIT[2346*9+8], INIT[2345*9+8], INIT[2344*9+8], 
           INIT[2343*9+8], INIT[2342*9+8], INIT[2341*9+8], INIT[2340*9+8], 
           INIT[2339*9+8], INIT[2338*9+8], INIT[2337*9+8], INIT[2336*9+8], 
           INIT[2335*9+8], INIT[2334*9+8], INIT[2333*9+8], INIT[2332*9+8], 
           INIT[2331*9+8], INIT[2330*9+8], INIT[2329*9+8], INIT[2328*9+8], 
           INIT[2327*9+8], INIT[2326*9+8], INIT[2325*9+8], INIT[2324*9+8], 
           INIT[2323*9+8], INIT[2322*9+8], INIT[2321*9+8], INIT[2320*9+8], 
           INIT[2319*9+8], INIT[2318*9+8], INIT[2317*9+8], INIT[2316*9+8], 
           INIT[2315*9+8], INIT[2314*9+8], INIT[2313*9+8], INIT[2312*9+8], 
           INIT[2311*9+8], INIT[2310*9+8], INIT[2309*9+8], INIT[2308*9+8], 
           INIT[2307*9+8], INIT[2306*9+8], INIT[2305*9+8], INIT[2304*9+8]}),
.INITP_0A({INIT[2815*9+8], INIT[2814*9+8], INIT[2813*9+8], INIT[2812*9+8], 
           INIT[2811*9+8], INIT[2810*9+8], INIT[2809*9+8], INIT[2808*9+8], 
           INIT[2807*9+8], INIT[2806*9+8], INIT[2805*9+8], INIT[2804*9+8], 
           INIT[2803*9+8], INIT[2802*9+8], INIT[2801*9+8], INIT[2800*9+8], 
           INIT[2799*9+8], INIT[2798*9+8], INIT[2797*9+8], INIT[2796*9+8], 
           INIT[2795*9+8], INIT[2794*9+8], INIT[2793*9+8], INIT[2792*9+8], 
           INIT[2791*9+8], INIT[2790*9+8], INIT[2789*9+8], INIT[2788*9+8], 
           INIT[2787*9+8], INIT[2786*9+8], INIT[2785*9+8], INIT[2784*9+8], 
           INIT[2783*9+8], INIT[2782*9+8], INIT[2781*9+8], INIT[2780*9+8], 
           INIT[2779*9+8], INIT[2778*9+8], INIT[2777*9+8], INIT[2776*9+8], 
           INIT[2775*9+8], INIT[2774*9+8], INIT[2773*9+8], INIT[2772*9+8], 
           INIT[2771*9+8], INIT[2770*9+8], INIT[2769*9+8], INIT[2768*9+8], 
           INIT[2767*9+8], INIT[2766*9+8], INIT[2765*9+8], INIT[2764*9+8], 
           INIT[2763*9+8], INIT[2762*9+8], INIT[2761*9+8], INIT[2760*9+8], 
           INIT[2759*9+8], INIT[2758*9+8], INIT[2757*9+8], INIT[2756*9+8], 
           INIT[2755*9+8], INIT[2754*9+8], INIT[2753*9+8], INIT[2752*9+8], 
           INIT[2751*9+8], INIT[2750*9+8], INIT[2749*9+8], INIT[2748*9+8], 
           INIT[2747*9+8], INIT[2746*9+8], INIT[2745*9+8], INIT[2744*9+8], 
           INIT[2743*9+8], INIT[2742*9+8], INIT[2741*9+8], INIT[2740*9+8], 
           INIT[2739*9+8], INIT[2738*9+8], INIT[2737*9+8], INIT[2736*9+8], 
           INIT[2735*9+8], INIT[2734*9+8], INIT[2733*9+8], INIT[2732*9+8], 
           INIT[2731*9+8], INIT[2730*9+8], INIT[2729*9+8], INIT[2728*9+8], 
           INIT[2727*9+8], INIT[2726*9+8], INIT[2725*9+8], INIT[2724*9+8], 
           INIT[2723*9+8], INIT[2722*9+8], INIT[2721*9+8], INIT[2720*9+8], 
           INIT[2719*9+8], INIT[2718*9+8], INIT[2717*9+8], INIT[2716*9+8], 
           INIT[2715*9+8], INIT[2714*9+8], INIT[2713*9+8], INIT[2712*9+8], 
           INIT[2711*9+8], INIT[2710*9+8], INIT[2709*9+8], INIT[2708*9+8], 
           INIT[2707*9+8], INIT[2706*9+8], INIT[2705*9+8], INIT[2704*9+8], 
           INIT[2703*9+8], INIT[2702*9+8], INIT[2701*9+8], INIT[2700*9+8], 
           INIT[2699*9+8], INIT[2698*9+8], INIT[2697*9+8], INIT[2696*9+8], 
           INIT[2695*9+8], INIT[2694*9+8], INIT[2693*9+8], INIT[2692*9+8], 
           INIT[2691*9+8], INIT[2690*9+8], INIT[2689*9+8], INIT[2688*9+8], 
           INIT[2687*9+8], INIT[2686*9+8], INIT[2685*9+8], INIT[2684*9+8], 
           INIT[2683*9+8], INIT[2682*9+8], INIT[2681*9+8], INIT[2680*9+8], 
           INIT[2679*9+8], INIT[2678*9+8], INIT[2677*9+8], INIT[2676*9+8], 
           INIT[2675*9+8], INIT[2674*9+8], INIT[2673*9+8], INIT[2672*9+8], 
           INIT[2671*9+8], INIT[2670*9+8], INIT[2669*9+8], INIT[2668*9+8], 
           INIT[2667*9+8], INIT[2666*9+8], INIT[2665*9+8], INIT[2664*9+8], 
           INIT[2663*9+8], INIT[2662*9+8], INIT[2661*9+8], INIT[2660*9+8], 
           INIT[2659*9+8], INIT[2658*9+8], INIT[2657*9+8], INIT[2656*9+8], 
           INIT[2655*9+8], INIT[2654*9+8], INIT[2653*9+8], INIT[2652*9+8], 
           INIT[2651*9+8], INIT[2650*9+8], INIT[2649*9+8], INIT[2648*9+8], 
           INIT[2647*9+8], INIT[2646*9+8], INIT[2645*9+8], INIT[2644*9+8], 
           INIT[2643*9+8], INIT[2642*9+8], INIT[2641*9+8], INIT[2640*9+8], 
           INIT[2639*9+8], INIT[2638*9+8], INIT[2637*9+8], INIT[2636*9+8], 
           INIT[2635*9+8], INIT[2634*9+8], INIT[2633*9+8], INIT[2632*9+8], 
           INIT[2631*9+8], INIT[2630*9+8], INIT[2629*9+8], INIT[2628*9+8], 
           INIT[2627*9+8], INIT[2626*9+8], INIT[2625*9+8], INIT[2624*9+8], 
           INIT[2623*9+8], INIT[2622*9+8], INIT[2621*9+8], INIT[2620*9+8], 
           INIT[2619*9+8], INIT[2618*9+8], INIT[2617*9+8], INIT[2616*9+8], 
           INIT[2615*9+8], INIT[2614*9+8], INIT[2613*9+8], INIT[2612*9+8], 
           INIT[2611*9+8], INIT[2610*9+8], INIT[2609*9+8], INIT[2608*9+8], 
           INIT[2607*9+8], INIT[2606*9+8], INIT[2605*9+8], INIT[2604*9+8], 
           INIT[2603*9+8], INIT[2602*9+8], INIT[2601*9+8], INIT[2600*9+8], 
           INIT[2599*9+8], INIT[2598*9+8], INIT[2597*9+8], INIT[2596*9+8], 
           INIT[2595*9+8], INIT[2594*9+8], INIT[2593*9+8], INIT[2592*9+8], 
           INIT[2591*9+8], INIT[2590*9+8], INIT[2589*9+8], INIT[2588*9+8], 
           INIT[2587*9+8], INIT[2586*9+8], INIT[2585*9+8], INIT[2584*9+8], 
           INIT[2583*9+8], INIT[2582*9+8], INIT[2581*9+8], INIT[2580*9+8], 
           INIT[2579*9+8], INIT[2578*9+8], INIT[2577*9+8], INIT[2576*9+8], 
           INIT[2575*9+8], INIT[2574*9+8], INIT[2573*9+8], INIT[2572*9+8], 
           INIT[2571*9+8], INIT[2570*9+8], INIT[2569*9+8], INIT[2568*9+8], 
           INIT[2567*9+8], INIT[2566*9+8], INIT[2565*9+8], INIT[2564*9+8], 
           INIT[2563*9+8], INIT[2562*9+8], INIT[2561*9+8], INIT[2560*9+8]}),
.INITP_0B({INIT[3071*9+8], INIT[3070*9+8], INIT[3069*9+8], INIT[3068*9+8], 
           INIT[3067*9+8], INIT[3066*9+8], INIT[3065*9+8], INIT[3064*9+8], 
           INIT[3063*9+8], INIT[3062*9+8], INIT[3061*9+8], INIT[3060*9+8], 
           INIT[3059*9+8], INIT[3058*9+8], INIT[3057*9+8], INIT[3056*9+8], 
           INIT[3055*9+8], INIT[3054*9+8], INIT[3053*9+8], INIT[3052*9+8], 
           INIT[3051*9+8], INIT[3050*9+8], INIT[3049*9+8], INIT[3048*9+8], 
           INIT[3047*9+8], INIT[3046*9+8], INIT[3045*9+8], INIT[3044*9+8], 
           INIT[3043*9+8], INIT[3042*9+8], INIT[3041*9+8], INIT[3040*9+8], 
           INIT[3039*9+8], INIT[3038*9+8], INIT[3037*9+8], INIT[3036*9+8], 
           INIT[3035*9+8], INIT[3034*9+8], INIT[3033*9+8], INIT[3032*9+8], 
           INIT[3031*9+8], INIT[3030*9+8], INIT[3029*9+8], INIT[3028*9+8], 
           INIT[3027*9+8], INIT[3026*9+8], INIT[3025*9+8], INIT[3024*9+8], 
           INIT[3023*9+8], INIT[3022*9+8], INIT[3021*9+8], INIT[3020*9+8], 
           INIT[3019*9+8], INIT[3018*9+8], INIT[3017*9+8], INIT[3016*9+8], 
           INIT[3015*9+8], INIT[3014*9+8], INIT[3013*9+8], INIT[3012*9+8], 
           INIT[3011*9+8], INIT[3010*9+8], INIT[3009*9+8], INIT[3008*9+8], 
           INIT[3007*9+8], INIT[3006*9+8], INIT[3005*9+8], INIT[3004*9+8], 
           INIT[3003*9+8], INIT[3002*9+8], INIT[3001*9+8], INIT[3000*9+8], 
           INIT[2999*9+8], INIT[2998*9+8], INIT[2997*9+8], INIT[2996*9+8], 
           INIT[2995*9+8], INIT[2994*9+8], INIT[2993*9+8], INIT[2992*9+8], 
           INIT[2991*9+8], INIT[2990*9+8], INIT[2989*9+8], INIT[2988*9+8], 
           INIT[2987*9+8], INIT[2986*9+8], INIT[2985*9+8], INIT[2984*9+8], 
           INIT[2983*9+8], INIT[2982*9+8], INIT[2981*9+8], INIT[2980*9+8], 
           INIT[2979*9+8], INIT[2978*9+8], INIT[2977*9+8], INIT[2976*9+8], 
           INIT[2975*9+8], INIT[2974*9+8], INIT[2973*9+8], INIT[2972*9+8], 
           INIT[2971*9+8], INIT[2970*9+8], INIT[2969*9+8], INIT[2968*9+8], 
           INIT[2967*9+8], INIT[2966*9+8], INIT[2965*9+8], INIT[2964*9+8], 
           INIT[2963*9+8], INIT[2962*9+8], INIT[2961*9+8], INIT[2960*9+8], 
           INIT[2959*9+8], INIT[2958*9+8], INIT[2957*9+8], INIT[2956*9+8], 
           INIT[2955*9+8], INIT[2954*9+8], INIT[2953*9+8], INIT[2952*9+8], 
           INIT[2951*9+8], INIT[2950*9+8], INIT[2949*9+8], INIT[2948*9+8], 
           INIT[2947*9+8], INIT[2946*9+8], INIT[2945*9+8], INIT[2944*9+8], 
           INIT[2943*9+8], INIT[2942*9+8], INIT[2941*9+8], INIT[2940*9+8], 
           INIT[2939*9+8], INIT[2938*9+8], INIT[2937*9+8], INIT[2936*9+8], 
           INIT[2935*9+8], INIT[2934*9+8], INIT[2933*9+8], INIT[2932*9+8], 
           INIT[2931*9+8], INIT[2930*9+8], INIT[2929*9+8], INIT[2928*9+8], 
           INIT[2927*9+8], INIT[2926*9+8], INIT[2925*9+8], INIT[2924*9+8], 
           INIT[2923*9+8], INIT[2922*9+8], INIT[2921*9+8], INIT[2920*9+8], 
           INIT[2919*9+8], INIT[2918*9+8], INIT[2917*9+8], INIT[2916*9+8], 
           INIT[2915*9+8], INIT[2914*9+8], INIT[2913*9+8], INIT[2912*9+8], 
           INIT[2911*9+8], INIT[2910*9+8], INIT[2909*9+8], INIT[2908*9+8], 
           INIT[2907*9+8], INIT[2906*9+8], INIT[2905*9+8], INIT[2904*9+8], 
           INIT[2903*9+8], INIT[2902*9+8], INIT[2901*9+8], INIT[2900*9+8], 
           INIT[2899*9+8], INIT[2898*9+8], INIT[2897*9+8], INIT[2896*9+8], 
           INIT[2895*9+8], INIT[2894*9+8], INIT[2893*9+8], INIT[2892*9+8], 
           INIT[2891*9+8], INIT[2890*9+8], INIT[2889*9+8], INIT[2888*9+8], 
           INIT[2887*9+8], INIT[2886*9+8], INIT[2885*9+8], INIT[2884*9+8], 
           INIT[2883*9+8], INIT[2882*9+8], INIT[2881*9+8], INIT[2880*9+8], 
           INIT[2879*9+8], INIT[2878*9+8], INIT[2877*9+8], INIT[2876*9+8], 
           INIT[2875*9+8], INIT[2874*9+8], INIT[2873*9+8], INIT[2872*9+8], 
           INIT[2871*9+8], INIT[2870*9+8], INIT[2869*9+8], INIT[2868*9+8], 
           INIT[2867*9+8], INIT[2866*9+8], INIT[2865*9+8], INIT[2864*9+8], 
           INIT[2863*9+8], INIT[2862*9+8], INIT[2861*9+8], INIT[2860*9+8], 
           INIT[2859*9+8], INIT[2858*9+8], INIT[2857*9+8], INIT[2856*9+8], 
           INIT[2855*9+8], INIT[2854*9+8], INIT[2853*9+8], INIT[2852*9+8], 
           INIT[2851*9+8], INIT[2850*9+8], INIT[2849*9+8], INIT[2848*9+8], 
           INIT[2847*9+8], INIT[2846*9+8], INIT[2845*9+8], INIT[2844*9+8], 
           INIT[2843*9+8], INIT[2842*9+8], INIT[2841*9+8], INIT[2840*9+8], 
           INIT[2839*9+8], INIT[2838*9+8], INIT[2837*9+8], INIT[2836*9+8], 
           INIT[2835*9+8], INIT[2834*9+8], INIT[2833*9+8], INIT[2832*9+8], 
           INIT[2831*9+8], INIT[2830*9+8], INIT[2829*9+8], INIT[2828*9+8], 
           INIT[2827*9+8], INIT[2826*9+8], INIT[2825*9+8], INIT[2824*9+8], 
           INIT[2823*9+8], INIT[2822*9+8], INIT[2821*9+8], INIT[2820*9+8], 
           INIT[2819*9+8], INIT[2818*9+8], INIT[2817*9+8], INIT[2816*9+8]}),
.INITP_0C({INIT[3327*9+8], INIT[3326*9+8], INIT[3325*9+8], INIT[3324*9+8], 
           INIT[3323*9+8], INIT[3322*9+8], INIT[3321*9+8], INIT[3320*9+8], 
           INIT[3319*9+8], INIT[3318*9+8], INIT[3317*9+8], INIT[3316*9+8], 
           INIT[3315*9+8], INIT[3314*9+8], INIT[3313*9+8], INIT[3312*9+8], 
           INIT[3311*9+8], INIT[3310*9+8], INIT[3309*9+8], INIT[3308*9+8], 
           INIT[3307*9+8], INIT[3306*9+8], INIT[3305*9+8], INIT[3304*9+8], 
           INIT[3303*9+8], INIT[3302*9+8], INIT[3301*9+8], INIT[3300*9+8], 
           INIT[3299*9+8], INIT[3298*9+8], INIT[3297*9+8], INIT[3296*9+8], 
           INIT[3295*9+8], INIT[3294*9+8], INIT[3293*9+8], INIT[3292*9+8], 
           INIT[3291*9+8], INIT[3290*9+8], INIT[3289*9+8], INIT[3288*9+8], 
           INIT[3287*9+8], INIT[3286*9+8], INIT[3285*9+8], INIT[3284*9+8], 
           INIT[3283*9+8], INIT[3282*9+8], INIT[3281*9+8], INIT[3280*9+8], 
           INIT[3279*9+8], INIT[3278*9+8], INIT[3277*9+8], INIT[3276*9+8], 
           INIT[3275*9+8], INIT[3274*9+8], INIT[3273*9+8], INIT[3272*9+8], 
           INIT[3271*9+8], INIT[3270*9+8], INIT[3269*9+8], INIT[3268*9+8], 
           INIT[3267*9+8], INIT[3266*9+8], INIT[3265*9+8], INIT[3264*9+8], 
           INIT[3263*9+8], INIT[3262*9+8], INIT[3261*9+8], INIT[3260*9+8], 
           INIT[3259*9+8], INIT[3258*9+8], INIT[3257*9+8], INIT[3256*9+8], 
           INIT[3255*9+8], INIT[3254*9+8], INIT[3253*9+8], INIT[3252*9+8], 
           INIT[3251*9+8], INIT[3250*9+8], INIT[3249*9+8], INIT[3248*9+8], 
           INIT[3247*9+8], INIT[3246*9+8], INIT[3245*9+8], INIT[3244*9+8], 
           INIT[3243*9+8], INIT[3242*9+8], INIT[3241*9+8], INIT[3240*9+8], 
           INIT[3239*9+8], INIT[3238*9+8], INIT[3237*9+8], INIT[3236*9+8], 
           INIT[3235*9+8], INIT[3234*9+8], INIT[3233*9+8], INIT[3232*9+8], 
           INIT[3231*9+8], INIT[3230*9+8], INIT[3229*9+8], INIT[3228*9+8], 
           INIT[3227*9+8], INIT[3226*9+8], INIT[3225*9+8], INIT[3224*9+8], 
           INIT[3223*9+8], INIT[3222*9+8], INIT[3221*9+8], INIT[3220*9+8], 
           INIT[3219*9+8], INIT[3218*9+8], INIT[3217*9+8], INIT[3216*9+8], 
           INIT[3215*9+8], INIT[3214*9+8], INIT[3213*9+8], INIT[3212*9+8], 
           INIT[3211*9+8], INIT[3210*9+8], INIT[3209*9+8], INIT[3208*9+8], 
           INIT[3207*9+8], INIT[3206*9+8], INIT[3205*9+8], INIT[3204*9+8], 
           INIT[3203*9+8], INIT[3202*9+8], INIT[3201*9+8], INIT[3200*9+8], 
           INIT[3199*9+8], INIT[3198*9+8], INIT[3197*9+8], INIT[3196*9+8], 
           INIT[3195*9+8], INIT[3194*9+8], INIT[3193*9+8], INIT[3192*9+8], 
           INIT[3191*9+8], INIT[3190*9+8], INIT[3189*9+8], INIT[3188*9+8], 
           INIT[3187*9+8], INIT[3186*9+8], INIT[3185*9+8], INIT[3184*9+8], 
           INIT[3183*9+8], INIT[3182*9+8], INIT[3181*9+8], INIT[3180*9+8], 
           INIT[3179*9+8], INIT[3178*9+8], INIT[3177*9+8], INIT[3176*9+8], 
           INIT[3175*9+8], INIT[3174*9+8], INIT[3173*9+8], INIT[3172*9+8], 
           INIT[3171*9+8], INIT[3170*9+8], INIT[3169*9+8], INIT[3168*9+8], 
           INIT[3167*9+8], INIT[3166*9+8], INIT[3165*9+8], INIT[3164*9+8], 
           INIT[3163*9+8], INIT[3162*9+8], INIT[3161*9+8], INIT[3160*9+8], 
           INIT[3159*9+8], INIT[3158*9+8], INIT[3157*9+8], INIT[3156*9+8], 
           INIT[3155*9+8], INIT[3154*9+8], INIT[3153*9+8], INIT[3152*9+8], 
           INIT[3151*9+8], INIT[3150*9+8], INIT[3149*9+8], INIT[3148*9+8], 
           INIT[3147*9+8], INIT[3146*9+8], INIT[3145*9+8], INIT[3144*9+8], 
           INIT[3143*9+8], INIT[3142*9+8], INIT[3141*9+8], INIT[3140*9+8], 
           INIT[3139*9+8], INIT[3138*9+8], INIT[3137*9+8], INIT[3136*9+8], 
           INIT[3135*9+8], INIT[3134*9+8], INIT[3133*9+8], INIT[3132*9+8], 
           INIT[3131*9+8], INIT[3130*9+8], INIT[3129*9+8], INIT[3128*9+8], 
           INIT[3127*9+8], INIT[3126*9+8], INIT[3125*9+8], INIT[3124*9+8], 
           INIT[3123*9+8], INIT[3122*9+8], INIT[3121*9+8], INIT[3120*9+8], 
           INIT[3119*9+8], INIT[3118*9+8], INIT[3117*9+8], INIT[3116*9+8], 
           INIT[3115*9+8], INIT[3114*9+8], INIT[3113*9+8], INIT[3112*9+8], 
           INIT[3111*9+8], INIT[3110*9+8], INIT[3109*9+8], INIT[3108*9+8], 
           INIT[3107*9+8], INIT[3106*9+8], INIT[3105*9+8], INIT[3104*9+8], 
           INIT[3103*9+8], INIT[3102*9+8], INIT[3101*9+8], INIT[3100*9+8], 
           INIT[3099*9+8], INIT[3098*9+8], INIT[3097*9+8], INIT[3096*9+8], 
           INIT[3095*9+8], INIT[3094*9+8], INIT[3093*9+8], INIT[3092*9+8], 
           INIT[3091*9+8], INIT[3090*9+8], INIT[3089*9+8], INIT[3088*9+8], 
           INIT[3087*9+8], INIT[3086*9+8], INIT[3085*9+8], INIT[3084*9+8], 
           INIT[3083*9+8], INIT[3082*9+8], INIT[3081*9+8], INIT[3080*9+8], 
           INIT[3079*9+8], INIT[3078*9+8], INIT[3077*9+8], INIT[3076*9+8], 
           INIT[3075*9+8], INIT[3074*9+8], INIT[3073*9+8], INIT[3072*9+8]}),
.INITP_0D({INIT[3583*9+8], INIT[3582*9+8], INIT[3581*9+8], INIT[3580*9+8], 
           INIT[3579*9+8], INIT[3578*9+8], INIT[3577*9+8], INIT[3576*9+8], 
           INIT[3575*9+8], INIT[3574*9+8], INIT[3573*9+8], INIT[3572*9+8], 
           INIT[3571*9+8], INIT[3570*9+8], INIT[3569*9+8], INIT[3568*9+8], 
           INIT[3567*9+8], INIT[3566*9+8], INIT[3565*9+8], INIT[3564*9+8], 
           INIT[3563*9+8], INIT[3562*9+8], INIT[3561*9+8], INIT[3560*9+8], 
           INIT[3559*9+8], INIT[3558*9+8], INIT[3557*9+8], INIT[3556*9+8], 
           INIT[3555*9+8], INIT[3554*9+8], INIT[3553*9+8], INIT[3552*9+8], 
           INIT[3551*9+8], INIT[3550*9+8], INIT[3549*9+8], INIT[3548*9+8], 
           INIT[3547*9+8], INIT[3546*9+8], INIT[3545*9+8], INIT[3544*9+8], 
           INIT[3543*9+8], INIT[3542*9+8], INIT[3541*9+8], INIT[3540*9+8], 
           INIT[3539*9+8], INIT[3538*9+8], INIT[3537*9+8], INIT[3536*9+8], 
           INIT[3535*9+8], INIT[3534*9+8], INIT[3533*9+8], INIT[3532*9+8], 
           INIT[3531*9+8], INIT[3530*9+8], INIT[3529*9+8], INIT[3528*9+8], 
           INIT[3527*9+8], INIT[3526*9+8], INIT[3525*9+8], INIT[3524*9+8], 
           INIT[3523*9+8], INIT[3522*9+8], INIT[3521*9+8], INIT[3520*9+8], 
           INIT[3519*9+8], INIT[3518*9+8], INIT[3517*9+8], INIT[3516*9+8], 
           INIT[3515*9+8], INIT[3514*9+8], INIT[3513*9+8], INIT[3512*9+8], 
           INIT[3511*9+8], INIT[3510*9+8], INIT[3509*9+8], INIT[3508*9+8], 
           INIT[3507*9+8], INIT[3506*9+8], INIT[3505*9+8], INIT[3504*9+8], 
           INIT[3503*9+8], INIT[3502*9+8], INIT[3501*9+8], INIT[3500*9+8], 
           INIT[3499*9+8], INIT[3498*9+8], INIT[3497*9+8], INIT[3496*9+8], 
           INIT[3495*9+8], INIT[3494*9+8], INIT[3493*9+8], INIT[3492*9+8], 
           INIT[3491*9+8], INIT[3490*9+8], INIT[3489*9+8], INIT[3488*9+8], 
           INIT[3487*9+8], INIT[3486*9+8], INIT[3485*9+8], INIT[3484*9+8], 
           INIT[3483*9+8], INIT[3482*9+8], INIT[3481*9+8], INIT[3480*9+8], 
           INIT[3479*9+8], INIT[3478*9+8], INIT[3477*9+8], INIT[3476*9+8], 
           INIT[3475*9+8], INIT[3474*9+8], INIT[3473*9+8], INIT[3472*9+8], 
           INIT[3471*9+8], INIT[3470*9+8], INIT[3469*9+8], INIT[3468*9+8], 
           INIT[3467*9+8], INIT[3466*9+8], INIT[3465*9+8], INIT[3464*9+8], 
           INIT[3463*9+8], INIT[3462*9+8], INIT[3461*9+8], INIT[3460*9+8], 
           INIT[3459*9+8], INIT[3458*9+8], INIT[3457*9+8], INIT[3456*9+8], 
           INIT[3455*9+8], INIT[3454*9+8], INIT[3453*9+8], INIT[3452*9+8], 
           INIT[3451*9+8], INIT[3450*9+8], INIT[3449*9+8], INIT[3448*9+8], 
           INIT[3447*9+8], INIT[3446*9+8], INIT[3445*9+8], INIT[3444*9+8], 
           INIT[3443*9+8], INIT[3442*9+8], INIT[3441*9+8], INIT[3440*9+8], 
           INIT[3439*9+8], INIT[3438*9+8], INIT[3437*9+8], INIT[3436*9+8], 
           INIT[3435*9+8], INIT[3434*9+8], INIT[3433*9+8], INIT[3432*9+8], 
           INIT[3431*9+8], INIT[3430*9+8], INIT[3429*9+8], INIT[3428*9+8], 
           INIT[3427*9+8], INIT[3426*9+8], INIT[3425*9+8], INIT[3424*9+8], 
           INIT[3423*9+8], INIT[3422*9+8], INIT[3421*9+8], INIT[3420*9+8], 
           INIT[3419*9+8], INIT[3418*9+8], INIT[3417*9+8], INIT[3416*9+8], 
           INIT[3415*9+8], INIT[3414*9+8], INIT[3413*9+8], INIT[3412*9+8], 
           INIT[3411*9+8], INIT[3410*9+8], INIT[3409*9+8], INIT[3408*9+8], 
           INIT[3407*9+8], INIT[3406*9+8], INIT[3405*9+8], INIT[3404*9+8], 
           INIT[3403*9+8], INIT[3402*9+8], INIT[3401*9+8], INIT[3400*9+8], 
           INIT[3399*9+8], INIT[3398*9+8], INIT[3397*9+8], INIT[3396*9+8], 
           INIT[3395*9+8], INIT[3394*9+8], INIT[3393*9+8], INIT[3392*9+8], 
           INIT[3391*9+8], INIT[3390*9+8], INIT[3389*9+8], INIT[3388*9+8], 
           INIT[3387*9+8], INIT[3386*9+8], INIT[3385*9+8], INIT[3384*9+8], 
           INIT[3383*9+8], INIT[3382*9+8], INIT[3381*9+8], INIT[3380*9+8], 
           INIT[3379*9+8], INIT[3378*9+8], INIT[3377*9+8], INIT[3376*9+8], 
           INIT[3375*9+8], INIT[3374*9+8], INIT[3373*9+8], INIT[3372*9+8], 
           INIT[3371*9+8], INIT[3370*9+8], INIT[3369*9+8], INIT[3368*9+8], 
           INIT[3367*9+8], INIT[3366*9+8], INIT[3365*9+8], INIT[3364*9+8], 
           INIT[3363*9+8], INIT[3362*9+8], INIT[3361*9+8], INIT[3360*9+8], 
           INIT[3359*9+8], INIT[3358*9+8], INIT[3357*9+8], INIT[3356*9+8], 
           INIT[3355*9+8], INIT[3354*9+8], INIT[3353*9+8], INIT[3352*9+8], 
           INIT[3351*9+8], INIT[3350*9+8], INIT[3349*9+8], INIT[3348*9+8], 
           INIT[3347*9+8], INIT[3346*9+8], INIT[3345*9+8], INIT[3344*9+8], 
           INIT[3343*9+8], INIT[3342*9+8], INIT[3341*9+8], INIT[3340*9+8], 
           INIT[3339*9+8], INIT[3338*9+8], INIT[3337*9+8], INIT[3336*9+8], 
           INIT[3335*9+8], INIT[3334*9+8], INIT[3333*9+8], INIT[3332*9+8], 
           INIT[3331*9+8], INIT[3330*9+8], INIT[3329*9+8], INIT[3328*9+8]}),
.INITP_0E({INIT[3839*9+8], INIT[3838*9+8], INIT[3837*9+8], INIT[3836*9+8], 
           INIT[3835*9+8], INIT[3834*9+8], INIT[3833*9+8], INIT[3832*9+8], 
           INIT[3831*9+8], INIT[3830*9+8], INIT[3829*9+8], INIT[3828*9+8], 
           INIT[3827*9+8], INIT[3826*9+8], INIT[3825*9+8], INIT[3824*9+8], 
           INIT[3823*9+8], INIT[3822*9+8], INIT[3821*9+8], INIT[3820*9+8], 
           INIT[3819*9+8], INIT[3818*9+8], INIT[3817*9+8], INIT[3816*9+8], 
           INIT[3815*9+8], INIT[3814*9+8], INIT[3813*9+8], INIT[3812*9+8], 
           INIT[3811*9+8], INIT[3810*9+8], INIT[3809*9+8], INIT[3808*9+8], 
           INIT[3807*9+8], INIT[3806*9+8], INIT[3805*9+8], INIT[3804*9+8], 
           INIT[3803*9+8], INIT[3802*9+8], INIT[3801*9+8], INIT[3800*9+8], 
           INIT[3799*9+8], INIT[3798*9+8], INIT[3797*9+8], INIT[3796*9+8], 
           INIT[3795*9+8], INIT[3794*9+8], INIT[3793*9+8], INIT[3792*9+8], 
           INIT[3791*9+8], INIT[3790*9+8], INIT[3789*9+8], INIT[3788*9+8], 
           INIT[3787*9+8], INIT[3786*9+8], INIT[3785*9+8], INIT[3784*9+8], 
           INIT[3783*9+8], INIT[3782*9+8], INIT[3781*9+8], INIT[3780*9+8], 
           INIT[3779*9+8], INIT[3778*9+8], INIT[3777*9+8], INIT[3776*9+8], 
           INIT[3775*9+8], INIT[3774*9+8], INIT[3773*9+8], INIT[3772*9+8], 
           INIT[3771*9+8], INIT[3770*9+8], INIT[3769*9+8], INIT[3768*9+8], 
           INIT[3767*9+8], INIT[3766*9+8], INIT[3765*9+8], INIT[3764*9+8], 
           INIT[3763*9+8], INIT[3762*9+8], INIT[3761*9+8], INIT[3760*9+8], 
           INIT[3759*9+8], INIT[3758*9+8], INIT[3757*9+8], INIT[3756*9+8], 
           INIT[3755*9+8], INIT[3754*9+8], INIT[3753*9+8], INIT[3752*9+8], 
           INIT[3751*9+8], INIT[3750*9+8], INIT[3749*9+8], INIT[3748*9+8], 
           INIT[3747*9+8], INIT[3746*9+8], INIT[3745*9+8], INIT[3744*9+8], 
           INIT[3743*9+8], INIT[3742*9+8], INIT[3741*9+8], INIT[3740*9+8], 
           INIT[3739*9+8], INIT[3738*9+8], INIT[3737*9+8], INIT[3736*9+8], 
           INIT[3735*9+8], INIT[3734*9+8], INIT[3733*9+8], INIT[3732*9+8], 
           INIT[3731*9+8], INIT[3730*9+8], INIT[3729*9+8], INIT[3728*9+8], 
           INIT[3727*9+8], INIT[3726*9+8], INIT[3725*9+8], INIT[3724*9+8], 
           INIT[3723*9+8], INIT[3722*9+8], INIT[3721*9+8], INIT[3720*9+8], 
           INIT[3719*9+8], INIT[3718*9+8], INIT[3717*9+8], INIT[3716*9+8], 
           INIT[3715*9+8], INIT[3714*9+8], INIT[3713*9+8], INIT[3712*9+8], 
           INIT[3711*9+8], INIT[3710*9+8], INIT[3709*9+8], INIT[3708*9+8], 
           INIT[3707*9+8], INIT[3706*9+8], INIT[3705*9+8], INIT[3704*9+8], 
           INIT[3703*9+8], INIT[3702*9+8], INIT[3701*9+8], INIT[3700*9+8], 
           INIT[3699*9+8], INIT[3698*9+8], INIT[3697*9+8], INIT[3696*9+8], 
           INIT[3695*9+8], INIT[3694*9+8], INIT[3693*9+8], INIT[3692*9+8], 
           INIT[3691*9+8], INIT[3690*9+8], INIT[3689*9+8], INIT[3688*9+8], 
           INIT[3687*9+8], INIT[3686*9+8], INIT[3685*9+8], INIT[3684*9+8], 
           INIT[3683*9+8], INIT[3682*9+8], INIT[3681*9+8], INIT[3680*9+8], 
           INIT[3679*9+8], INIT[3678*9+8], INIT[3677*9+8], INIT[3676*9+8], 
           INIT[3675*9+8], INIT[3674*9+8], INIT[3673*9+8], INIT[3672*9+8], 
           INIT[3671*9+8], INIT[3670*9+8], INIT[3669*9+8], INIT[3668*9+8], 
           INIT[3667*9+8], INIT[3666*9+8], INIT[3665*9+8], INIT[3664*9+8], 
           INIT[3663*9+8], INIT[3662*9+8], INIT[3661*9+8], INIT[3660*9+8], 
           INIT[3659*9+8], INIT[3658*9+8], INIT[3657*9+8], INIT[3656*9+8], 
           INIT[3655*9+8], INIT[3654*9+8], INIT[3653*9+8], INIT[3652*9+8], 
           INIT[3651*9+8], INIT[3650*9+8], INIT[3649*9+8], INIT[3648*9+8], 
           INIT[3647*9+8], INIT[3646*9+8], INIT[3645*9+8], INIT[3644*9+8], 
           INIT[3643*9+8], INIT[3642*9+8], INIT[3641*9+8], INIT[3640*9+8], 
           INIT[3639*9+8], INIT[3638*9+8], INIT[3637*9+8], INIT[3636*9+8], 
           INIT[3635*9+8], INIT[3634*9+8], INIT[3633*9+8], INIT[3632*9+8], 
           INIT[3631*9+8], INIT[3630*9+8], INIT[3629*9+8], INIT[3628*9+8], 
           INIT[3627*9+8], INIT[3626*9+8], INIT[3625*9+8], INIT[3624*9+8], 
           INIT[3623*9+8], INIT[3622*9+8], INIT[3621*9+8], INIT[3620*9+8], 
           INIT[3619*9+8], INIT[3618*9+8], INIT[3617*9+8], INIT[3616*9+8], 
           INIT[3615*9+8], INIT[3614*9+8], INIT[3613*9+8], INIT[3612*9+8], 
           INIT[3611*9+8], INIT[3610*9+8], INIT[3609*9+8], INIT[3608*9+8], 
           INIT[3607*9+8], INIT[3606*9+8], INIT[3605*9+8], INIT[3604*9+8], 
           INIT[3603*9+8], INIT[3602*9+8], INIT[3601*9+8], INIT[3600*9+8], 
           INIT[3599*9+8], INIT[3598*9+8], INIT[3597*9+8], INIT[3596*9+8], 
           INIT[3595*9+8], INIT[3594*9+8], INIT[3593*9+8], INIT[3592*9+8], 
           INIT[3591*9+8], INIT[3590*9+8], INIT[3589*9+8], INIT[3588*9+8], 
           INIT[3587*9+8], INIT[3586*9+8], INIT[3585*9+8], INIT[3584*9+8]}),
.INITP_0F({INIT[4095*9+8], INIT[4094*9+8], INIT[4093*9+8], INIT[4092*9+8], 
           INIT[4091*9+8], INIT[4090*9+8], INIT[4089*9+8], INIT[4088*9+8], 
           INIT[4087*9+8], INIT[4086*9+8], INIT[4085*9+8], INIT[4084*9+8], 
           INIT[4083*9+8], INIT[4082*9+8], INIT[4081*9+8], INIT[4080*9+8], 
           INIT[4079*9+8], INIT[4078*9+8], INIT[4077*9+8], INIT[4076*9+8], 
           INIT[4075*9+8], INIT[4074*9+8], INIT[4073*9+8], INIT[4072*9+8], 
           INIT[4071*9+8], INIT[4070*9+8], INIT[4069*9+8], INIT[4068*9+8], 
           INIT[4067*9+8], INIT[4066*9+8], INIT[4065*9+8], INIT[4064*9+8], 
           INIT[4063*9+8], INIT[4062*9+8], INIT[4061*9+8], INIT[4060*9+8], 
           INIT[4059*9+8], INIT[4058*9+8], INIT[4057*9+8], INIT[4056*9+8], 
           INIT[4055*9+8], INIT[4054*9+8], INIT[4053*9+8], INIT[4052*9+8], 
           INIT[4051*9+8], INIT[4050*9+8], INIT[4049*9+8], INIT[4048*9+8], 
           INIT[4047*9+8], INIT[4046*9+8], INIT[4045*9+8], INIT[4044*9+8], 
           INIT[4043*9+8], INIT[4042*9+8], INIT[4041*9+8], INIT[4040*9+8], 
           INIT[4039*9+8], INIT[4038*9+8], INIT[4037*9+8], INIT[4036*9+8], 
           INIT[4035*9+8], INIT[4034*9+8], INIT[4033*9+8], INIT[4032*9+8], 
           INIT[4031*9+8], INIT[4030*9+8], INIT[4029*9+8], INIT[4028*9+8], 
           INIT[4027*9+8], INIT[4026*9+8], INIT[4025*9+8], INIT[4024*9+8], 
           INIT[4023*9+8], INIT[4022*9+8], INIT[4021*9+8], INIT[4020*9+8], 
           INIT[4019*9+8], INIT[4018*9+8], INIT[4017*9+8], INIT[4016*9+8], 
           INIT[4015*9+8], INIT[4014*9+8], INIT[4013*9+8], INIT[4012*9+8], 
           INIT[4011*9+8], INIT[4010*9+8], INIT[4009*9+8], INIT[4008*9+8], 
           INIT[4007*9+8], INIT[4006*9+8], INIT[4005*9+8], INIT[4004*9+8], 
           INIT[4003*9+8], INIT[4002*9+8], INIT[4001*9+8], INIT[4000*9+8], 
           INIT[3999*9+8], INIT[3998*9+8], INIT[3997*9+8], INIT[3996*9+8], 
           INIT[3995*9+8], INIT[3994*9+8], INIT[3993*9+8], INIT[3992*9+8], 
           INIT[3991*9+8], INIT[3990*9+8], INIT[3989*9+8], INIT[3988*9+8], 
           INIT[3987*9+8], INIT[3986*9+8], INIT[3985*9+8], INIT[3984*9+8], 
           INIT[3983*9+8], INIT[3982*9+8], INIT[3981*9+8], INIT[3980*9+8], 
           INIT[3979*9+8], INIT[3978*9+8], INIT[3977*9+8], INIT[3976*9+8], 
           INIT[3975*9+8], INIT[3974*9+8], INIT[3973*9+8], INIT[3972*9+8], 
           INIT[3971*9+8], INIT[3970*9+8], INIT[3969*9+8], INIT[3968*9+8], 
           INIT[3967*9+8], INIT[3966*9+8], INIT[3965*9+8], INIT[3964*9+8], 
           INIT[3963*9+8], INIT[3962*9+8], INIT[3961*9+8], INIT[3960*9+8], 
           INIT[3959*9+8], INIT[3958*9+8], INIT[3957*9+8], INIT[3956*9+8], 
           INIT[3955*9+8], INIT[3954*9+8], INIT[3953*9+8], INIT[3952*9+8], 
           INIT[3951*9+8], INIT[3950*9+8], INIT[3949*9+8], INIT[3948*9+8], 
           INIT[3947*9+8], INIT[3946*9+8], INIT[3945*9+8], INIT[3944*9+8], 
           INIT[3943*9+8], INIT[3942*9+8], INIT[3941*9+8], INIT[3940*9+8], 
           INIT[3939*9+8], INIT[3938*9+8], INIT[3937*9+8], INIT[3936*9+8], 
           INIT[3935*9+8], INIT[3934*9+8], INIT[3933*9+8], INIT[3932*9+8], 
           INIT[3931*9+8], INIT[3930*9+8], INIT[3929*9+8], INIT[3928*9+8], 
           INIT[3927*9+8], INIT[3926*9+8], INIT[3925*9+8], INIT[3924*9+8], 
           INIT[3923*9+8], INIT[3922*9+8], INIT[3921*9+8], INIT[3920*9+8], 
           INIT[3919*9+8], INIT[3918*9+8], INIT[3917*9+8], INIT[3916*9+8], 
           INIT[3915*9+8], INIT[3914*9+8], INIT[3913*9+8], INIT[3912*9+8], 
           INIT[3911*9+8], INIT[3910*9+8], INIT[3909*9+8], INIT[3908*9+8], 
           INIT[3907*9+8], INIT[3906*9+8], INIT[3905*9+8], INIT[3904*9+8], 
           INIT[3903*9+8], INIT[3902*9+8], INIT[3901*9+8], INIT[3900*9+8], 
           INIT[3899*9+8], INIT[3898*9+8], INIT[3897*9+8], INIT[3896*9+8], 
           INIT[3895*9+8], INIT[3894*9+8], INIT[3893*9+8], INIT[3892*9+8], 
           INIT[3891*9+8], INIT[3890*9+8], INIT[3889*9+8], INIT[3888*9+8], 
           INIT[3887*9+8], INIT[3886*9+8], INIT[3885*9+8], INIT[3884*9+8], 
           INIT[3883*9+8], INIT[3882*9+8], INIT[3881*9+8], INIT[3880*9+8], 
           INIT[3879*9+8], INIT[3878*9+8], INIT[3877*9+8], INIT[3876*9+8], 
           INIT[3875*9+8], INIT[3874*9+8], INIT[3873*9+8], INIT[3872*9+8], 
           INIT[3871*9+8], INIT[3870*9+8], INIT[3869*9+8], INIT[3868*9+8], 
           INIT[3867*9+8], INIT[3866*9+8], INIT[3865*9+8], INIT[3864*9+8], 
           INIT[3863*9+8], INIT[3862*9+8], INIT[3861*9+8], INIT[3860*9+8], 
           INIT[3859*9+8], INIT[3858*9+8], INIT[3857*9+8], INIT[3856*9+8], 
           INIT[3855*9+8], INIT[3854*9+8], INIT[3853*9+8], INIT[3852*9+8], 
           INIT[3851*9+8], INIT[3850*9+8], INIT[3849*9+8], INIT[3848*9+8], 
           INIT[3847*9+8], INIT[3846*9+8], INIT[3845*9+8], INIT[3844*9+8], 
           INIT[3843*9+8], INIT[3842*9+8], INIT[3841*9+8], INIT[3840*9+8]}),
.INIT_00({INIT[ 31*9 +: 8], INIT[ 30*9 +: 8], INIT[ 29*9 +: 8], INIT[ 28*9 +: 8], 
          INIT[ 27*9 +: 8], INIT[ 26*9 +: 8], INIT[ 25*9 +: 8], INIT[ 24*9 +: 8], 
          INIT[ 23*9 +: 8], INIT[ 22*9 +: 8], INIT[ 21*9 +: 8], INIT[ 20*9 +: 8], 
          INIT[ 19*9 +: 8], INIT[ 18*9 +: 8], INIT[ 17*9 +: 8], INIT[ 16*9 +: 8], 
          INIT[ 15*9 +: 8], INIT[ 14*9 +: 8], INIT[ 13*9 +: 8], INIT[ 12*9 +: 8], 
          INIT[ 11*9 +: 8], INIT[ 10*9 +: 8], INIT[  9*9 +: 8], INIT[  8*9 +: 8], 
          INIT[  7*9 +: 8], INIT[  6*9 +: 8], INIT[  5*9 +: 8], INIT[  4*9 +: 8], 
          INIT[  3*9 +: 8], INIT[  2*9 +: 8], INIT[  1*9 +: 8], INIT[  0*9 +: 8]}),
.INIT_01({INIT[ 63*9 +: 8], INIT[ 62*9 +: 8], INIT[ 61*9 +: 8], INIT[ 60*9 +: 8], 
          INIT[ 59*9 +: 8], INIT[ 58*9 +: 8], INIT[ 57*9 +: 8], INIT[ 56*9 +: 8], 
          INIT[ 55*9 +: 8], INIT[ 54*9 +: 8], INIT[ 53*9 +: 8], INIT[ 52*9 +: 8], 
          INIT[ 51*9 +: 8], INIT[ 50*9 +: 8], INIT[ 49*9 +: 8], INIT[ 48*9 +: 8], 
          INIT[ 47*9 +: 8], INIT[ 46*9 +: 8], INIT[ 45*9 +: 8], INIT[ 44*9 +: 8], 
          INIT[ 43*9 +: 8], INIT[ 42*9 +: 8], INIT[ 41*9 +: 8], INIT[ 40*9 +: 8], 
          INIT[ 39*9 +: 8], INIT[ 38*9 +: 8], INIT[ 37*9 +: 8], INIT[ 36*9 +: 8], 
          INIT[ 35*9 +: 8], INIT[ 34*9 +: 8], INIT[ 33*9 +: 8], INIT[ 32*9 +: 8]}),
.INIT_02({INIT[ 95*9 +: 8], INIT[ 94*9 +: 8], INIT[ 93*9 +: 8], INIT[ 92*9 +: 8], 
          INIT[ 91*9 +: 8], INIT[ 90*9 +: 8], INIT[ 89*9 +: 8], INIT[ 88*9 +: 8], 
          INIT[ 87*9 +: 8], INIT[ 86*9 +: 8], INIT[ 85*9 +: 8], INIT[ 84*9 +: 8], 
          INIT[ 83*9 +: 8], INIT[ 82*9 +: 8], INIT[ 81*9 +: 8], INIT[ 80*9 +: 8], 
          INIT[ 79*9 +: 8], INIT[ 78*9 +: 8], INIT[ 77*9 +: 8], INIT[ 76*9 +: 8], 
          INIT[ 75*9 +: 8], INIT[ 74*9 +: 8], INIT[ 73*9 +: 8], INIT[ 72*9 +: 8], 
          INIT[ 71*9 +: 8], INIT[ 70*9 +: 8], INIT[ 69*9 +: 8], INIT[ 68*9 +: 8], 
          INIT[ 67*9 +: 8], INIT[ 66*9 +: 8], INIT[ 65*9 +: 8], INIT[ 64*9 +: 8]}),
.INIT_03({INIT[127*9 +: 8], INIT[126*9 +: 8], INIT[125*9 +: 8], INIT[124*9 +: 8], 
          INIT[123*9 +: 8], INIT[122*9 +: 8], INIT[121*9 +: 8], INIT[120*9 +: 8], 
          INIT[119*9 +: 8], INIT[118*9 +: 8], INIT[117*9 +: 8], INIT[116*9 +: 8], 
          INIT[115*9 +: 8], INIT[114*9 +: 8], INIT[113*9 +: 8], INIT[112*9 +: 8], 
          INIT[111*9 +: 8], INIT[110*9 +: 8], INIT[109*9 +: 8], INIT[108*9 +: 8], 
          INIT[107*9 +: 8], INIT[106*9 +: 8], INIT[105*9 +: 8], INIT[104*9 +: 8], 
          INIT[103*9 +: 8], INIT[102*9 +: 8], INIT[101*9 +: 8], INIT[100*9 +: 8], 
          INIT[ 99*9 +: 8], INIT[ 98*9 +: 8], INIT[ 97*9 +: 8], INIT[ 96*9 +: 8]}),
.INIT_04({INIT[159*9 +: 8], INIT[158*9 +: 8], INIT[157*9 +: 8], INIT[156*9 +: 8], 
          INIT[155*9 +: 8], INIT[154*9 +: 8], INIT[153*9 +: 8], INIT[152*9 +: 8], 
          INIT[151*9 +: 8], INIT[150*9 +: 8], INIT[149*9 +: 8], INIT[148*9 +: 8], 
          INIT[147*9 +: 8], INIT[146*9 +: 8], INIT[145*9 +: 8], INIT[144*9 +: 8], 
          INIT[143*9 +: 8], INIT[142*9 +: 8], INIT[141*9 +: 8], INIT[140*9 +: 8], 
          INIT[139*9 +: 8], INIT[138*9 +: 8], INIT[137*9 +: 8], INIT[136*9 +: 8], 
          INIT[135*9 +: 8], INIT[134*9 +: 8], INIT[133*9 +: 8], INIT[132*9 +: 8], 
          INIT[131*9 +: 8], INIT[130*9 +: 8], INIT[129*9 +: 8], INIT[128*9 +: 8]}),
.INIT_05({INIT[191*9 +: 8], INIT[190*9 +: 8], INIT[189*9 +: 8], INIT[188*9 +: 8], 
          INIT[187*9 +: 8], INIT[186*9 +: 8], INIT[185*9 +: 8], INIT[184*9 +: 8], 
          INIT[183*9 +: 8], INIT[182*9 +: 8], INIT[181*9 +: 8], INIT[180*9 +: 8], 
          INIT[179*9 +: 8], INIT[178*9 +: 8], INIT[177*9 +: 8], INIT[176*9 +: 8], 
          INIT[175*9 +: 8], INIT[174*9 +: 8], INIT[173*9 +: 8], INIT[172*9 +: 8], 
          INIT[171*9 +: 8], INIT[170*9 +: 8], INIT[169*9 +: 8], INIT[168*9 +: 8], 
          INIT[167*9 +: 8], INIT[166*9 +: 8], INIT[165*9 +: 8], INIT[164*9 +: 8], 
          INIT[163*9 +: 8], INIT[162*9 +: 8], INIT[161*9 +: 8], INIT[160*9 +: 8]}),
.INIT_06({INIT[223*9 +: 8], INIT[222*9 +: 8], INIT[221*9 +: 8], INIT[220*9 +: 8], 
          INIT[219*9 +: 8], INIT[218*9 +: 8], INIT[217*9 +: 8], INIT[216*9 +: 8], 
          INIT[215*9 +: 8], INIT[214*9 +: 8], INIT[213*9 +: 8], INIT[212*9 +: 8], 
          INIT[211*9 +: 8], INIT[210*9 +: 8], INIT[209*9 +: 8], INIT[208*9 +: 8], 
          INIT[207*9 +: 8], INIT[206*9 +: 8], INIT[205*9 +: 8], INIT[204*9 +: 8], 
          INIT[203*9 +: 8], INIT[202*9 +: 8], INIT[201*9 +: 8], INIT[200*9 +: 8], 
          INIT[199*9 +: 8], INIT[198*9 +: 8], INIT[197*9 +: 8], INIT[196*9 +: 8], 
          INIT[195*9 +: 8], INIT[194*9 +: 8], INIT[193*9 +: 8], INIT[192*9 +: 8]}),
.INIT_07({INIT[255*9 +: 8], INIT[254*9 +: 8], INIT[253*9 +: 8], INIT[252*9 +: 8], 
          INIT[251*9 +: 8], INIT[250*9 +: 8], INIT[249*9 +: 8], INIT[248*9 +: 8], 
          INIT[247*9 +: 8], INIT[246*9 +: 8], INIT[245*9 +: 8], INIT[244*9 +: 8], 
          INIT[243*9 +: 8], INIT[242*9 +: 8], INIT[241*9 +: 8], INIT[240*9 +: 8], 
          INIT[239*9 +: 8], INIT[238*9 +: 8], INIT[237*9 +: 8], INIT[236*9 +: 8], 
          INIT[235*9 +: 8], INIT[234*9 +: 8], INIT[233*9 +: 8], INIT[232*9 +: 8], 
          INIT[231*9 +: 8], INIT[230*9 +: 8], INIT[229*9 +: 8], INIT[228*9 +: 8], 
          INIT[227*9 +: 8], INIT[226*9 +: 8], INIT[225*9 +: 8], INIT[224*9 +: 8]}),
.INIT_08({INIT[287*9 +: 8], INIT[286*9 +: 8], INIT[285*9 +: 8], INIT[284*9 +: 8], 
          INIT[283*9 +: 8], INIT[282*9 +: 8], INIT[281*9 +: 8], INIT[280*9 +: 8], 
          INIT[279*9 +: 8], INIT[278*9 +: 8], INIT[277*9 +: 8], INIT[276*9 +: 8], 
          INIT[275*9 +: 8], INIT[274*9 +: 8], INIT[273*9 +: 8], INIT[272*9 +: 8], 
          INIT[271*9 +: 8], INIT[270*9 +: 8], INIT[269*9 +: 8], INIT[268*9 +: 8], 
          INIT[267*9 +: 8], INIT[266*9 +: 8], INIT[265*9 +: 8], INIT[264*9 +: 8], 
          INIT[263*9 +: 8], INIT[262*9 +: 8], INIT[261*9 +: 8], INIT[260*9 +: 8], 
          INIT[259*9 +: 8], INIT[258*9 +: 8], INIT[257*9 +: 8], INIT[256*9 +: 8]}),
.INIT_09({INIT[319*9 +: 8], INIT[318*9 +: 8], INIT[317*9 +: 8], INIT[316*9 +: 8], 
          INIT[315*9 +: 8], INIT[314*9 +: 8], INIT[313*9 +: 8], INIT[312*9 +: 8], 
          INIT[311*9 +: 8], INIT[310*9 +: 8], INIT[309*9 +: 8], INIT[308*9 +: 8], 
          INIT[307*9 +: 8], INIT[306*9 +: 8], INIT[305*9 +: 8], INIT[304*9 +: 8], 
          INIT[303*9 +: 8], INIT[302*9 +: 8], INIT[301*9 +: 8], INIT[300*9 +: 8], 
          INIT[299*9 +: 8], INIT[298*9 +: 8], INIT[297*9 +: 8], INIT[296*9 +: 8], 
          INIT[295*9 +: 8], INIT[294*9 +: 8], INIT[293*9 +: 8], INIT[292*9 +: 8], 
          INIT[291*9 +: 8], INIT[290*9 +: 8], INIT[289*9 +: 8], INIT[288*9 +: 8]}),
.INIT_0A({INIT[351*9 +: 8], INIT[350*9 +: 8], INIT[349*9 +: 8], INIT[348*9 +: 8], 
          INIT[347*9 +: 8], INIT[346*9 +: 8], INIT[345*9 +: 8], INIT[344*9 +: 8], 
          INIT[343*9 +: 8], INIT[342*9 +: 8], INIT[341*9 +: 8], INIT[340*9 +: 8], 
          INIT[339*9 +: 8], INIT[338*9 +: 8], INIT[337*9 +: 8], INIT[336*9 +: 8], 
          INIT[335*9 +: 8], INIT[334*9 +: 8], INIT[333*9 +: 8], INIT[332*9 +: 8], 
          INIT[331*9 +: 8], INIT[330*9 +: 8], INIT[329*9 +: 8], INIT[328*9 +: 8], 
          INIT[327*9 +: 8], INIT[326*9 +: 8], INIT[325*9 +: 8], INIT[324*9 +: 8], 
          INIT[323*9 +: 8], INIT[322*9 +: 8], INIT[321*9 +: 8], INIT[320*9 +: 8]}),
.INIT_0B({INIT[383*9 +: 8], INIT[382*9 +: 8], INIT[381*9 +: 8], INIT[380*9 +: 8], 
          INIT[379*9 +: 8], INIT[378*9 +: 8], INIT[377*9 +: 8], INIT[376*9 +: 8], 
          INIT[375*9 +: 8], INIT[374*9 +: 8], INIT[373*9 +: 8], INIT[372*9 +: 8], 
          INIT[371*9 +: 8], INIT[370*9 +: 8], INIT[369*9 +: 8], INIT[368*9 +: 8], 
          INIT[367*9 +: 8], INIT[366*9 +: 8], INIT[365*9 +: 8], INIT[364*9 +: 8], 
          INIT[363*9 +: 8], INIT[362*9 +: 8], INIT[361*9 +: 8], INIT[360*9 +: 8], 
          INIT[359*9 +: 8], INIT[358*9 +: 8], INIT[357*9 +: 8], INIT[356*9 +: 8], 
          INIT[355*9 +: 8], INIT[354*9 +: 8], INIT[353*9 +: 8], INIT[352*9 +: 8]}),
.INIT_0C({INIT[415*9 +: 8], INIT[414*9 +: 8], INIT[413*9 +: 8], INIT[412*9 +: 8], 
          INIT[411*9 +: 8], INIT[410*9 +: 8], INIT[409*9 +: 8], INIT[408*9 +: 8], 
          INIT[407*9 +: 8], INIT[406*9 +: 8], INIT[405*9 +: 8], INIT[404*9 +: 8], 
          INIT[403*9 +: 8], INIT[402*9 +: 8], INIT[401*9 +: 8], INIT[400*9 +: 8], 
          INIT[399*9 +: 8], INIT[398*9 +: 8], INIT[397*9 +: 8], INIT[396*9 +: 8], 
          INIT[395*9 +: 8], INIT[394*9 +: 8], INIT[393*9 +: 8], INIT[392*9 +: 8], 
          INIT[391*9 +: 8], INIT[390*9 +: 8], INIT[389*9 +: 8], INIT[388*9 +: 8], 
          INIT[387*9 +: 8], INIT[386*9 +: 8], INIT[385*9 +: 8], INIT[384*9 +: 8]}),
.INIT_0D({INIT[447*9 +: 8], INIT[446*9 +: 8], INIT[445*9 +: 8], INIT[444*9 +: 8], 
          INIT[443*9 +: 8], INIT[442*9 +: 8], INIT[441*9 +: 8], INIT[440*9 +: 8], 
          INIT[439*9 +: 8], INIT[438*9 +: 8], INIT[437*9 +: 8], INIT[436*9 +: 8], 
          INIT[435*9 +: 8], INIT[434*9 +: 8], INIT[433*9 +: 8], INIT[432*9 +: 8], 
          INIT[431*9 +: 8], INIT[430*9 +: 8], INIT[429*9 +: 8], INIT[428*9 +: 8], 
          INIT[427*9 +: 8], INIT[426*9 +: 8], INIT[425*9 +: 8], INIT[424*9 +: 8], 
          INIT[423*9 +: 8], INIT[422*9 +: 8], INIT[421*9 +: 8], INIT[420*9 +: 8], 
          INIT[419*9 +: 8], INIT[418*9 +: 8], INIT[417*9 +: 8], INIT[416*9 +: 8]}),
.INIT_0E({INIT[479*9 +: 8], INIT[478*9 +: 8], INIT[477*9 +: 8], INIT[476*9 +: 8], 
          INIT[475*9 +: 8], INIT[474*9 +: 8], INIT[473*9 +: 8], INIT[472*9 +: 8], 
          INIT[471*9 +: 8], INIT[470*9 +: 8], INIT[469*9 +: 8], INIT[468*9 +: 8], 
          INIT[467*9 +: 8], INIT[466*9 +: 8], INIT[465*9 +: 8], INIT[464*9 +: 8], 
          INIT[463*9 +: 8], INIT[462*9 +: 8], INIT[461*9 +: 8], INIT[460*9 +: 8], 
          INIT[459*9 +: 8], INIT[458*9 +: 8], INIT[457*9 +: 8], INIT[456*9 +: 8], 
          INIT[455*9 +: 8], INIT[454*9 +: 8], INIT[453*9 +: 8], INIT[452*9 +: 8], 
          INIT[451*9 +: 8], INIT[450*9 +: 8], INIT[449*9 +: 8], INIT[448*9 +: 8]}),
.INIT_0F({INIT[511*9 +: 8], INIT[510*9 +: 8], INIT[509*9 +: 8], INIT[508*9 +: 8], 
          INIT[507*9 +: 8], INIT[506*9 +: 8], INIT[505*9 +: 8], INIT[504*9 +: 8], 
          INIT[503*9 +: 8], INIT[502*9 +: 8], INIT[501*9 +: 8], INIT[500*9 +: 8], 
          INIT[499*9 +: 8], INIT[498*9 +: 8], INIT[497*9 +: 8], INIT[496*9 +: 8], 
          INIT[495*9 +: 8], INIT[494*9 +: 8], INIT[493*9 +: 8], INIT[492*9 +: 8], 
          INIT[491*9 +: 8], INIT[490*9 +: 8], INIT[489*9 +: 8], INIT[488*9 +: 8], 
          INIT[487*9 +: 8], INIT[486*9 +: 8], INIT[485*9 +: 8], INIT[484*9 +: 8], 
          INIT[483*9 +: 8], INIT[482*9 +: 8], INIT[481*9 +: 8], INIT[480*9 +: 8]}),
.INIT_10({INIT[543*9 +: 8], INIT[542*9 +: 8], INIT[541*9 +: 8], INIT[540*9 +: 8], 
          INIT[539*9 +: 8], INIT[538*9 +: 8], INIT[537*9 +: 8], INIT[536*9 +: 8], 
          INIT[535*9 +: 8], INIT[534*9 +: 8], INIT[533*9 +: 8], INIT[532*9 +: 8], 
          INIT[531*9 +: 8], INIT[530*9 +: 8], INIT[529*9 +: 8], INIT[528*9 +: 8], 
          INIT[527*9 +: 8], INIT[526*9 +: 8], INIT[525*9 +: 8], INIT[524*9 +: 8], 
          INIT[523*9 +: 8], INIT[522*9 +: 8], INIT[521*9 +: 8], INIT[520*9 +: 8], 
          INIT[519*9 +: 8], INIT[518*9 +: 8], INIT[517*9 +: 8], INIT[516*9 +: 8], 
          INIT[515*9 +: 8], INIT[514*9 +: 8], INIT[513*9 +: 8], INIT[512*9 +: 8]}),
.INIT_11({INIT[575*9 +: 8], INIT[574*9 +: 8], INIT[573*9 +: 8], INIT[572*9 +: 8], 
          INIT[571*9 +: 8], INIT[570*9 +: 8], INIT[569*9 +: 8], INIT[568*9 +: 8], 
          INIT[567*9 +: 8], INIT[566*9 +: 8], INIT[565*9 +: 8], INIT[564*9 +: 8], 
          INIT[563*9 +: 8], INIT[562*9 +: 8], INIT[561*9 +: 8], INIT[560*9 +: 8], 
          INIT[559*9 +: 8], INIT[558*9 +: 8], INIT[557*9 +: 8], INIT[556*9 +: 8], 
          INIT[555*9 +: 8], INIT[554*9 +: 8], INIT[553*9 +: 8], INIT[552*9 +: 8], 
          INIT[551*9 +: 8], INIT[550*9 +: 8], INIT[549*9 +: 8], INIT[548*9 +: 8], 
          INIT[547*9 +: 8], INIT[546*9 +: 8], INIT[545*9 +: 8], INIT[544*9 +: 8]}),
.INIT_12({INIT[607*9 +: 8], INIT[606*9 +: 8], INIT[605*9 +: 8], INIT[604*9 +: 8], 
          INIT[603*9 +: 8], INIT[602*9 +: 8], INIT[601*9 +: 8], INIT[600*9 +: 8], 
          INIT[599*9 +: 8], INIT[598*9 +: 8], INIT[597*9 +: 8], INIT[596*9 +: 8], 
          INIT[595*9 +: 8], INIT[594*9 +: 8], INIT[593*9 +: 8], INIT[592*9 +: 8], 
          INIT[591*9 +: 8], INIT[590*9 +: 8], INIT[589*9 +: 8], INIT[588*9 +: 8], 
          INIT[587*9 +: 8], INIT[586*9 +: 8], INIT[585*9 +: 8], INIT[584*9 +: 8], 
          INIT[583*9 +: 8], INIT[582*9 +: 8], INIT[581*9 +: 8], INIT[580*9 +: 8], 
          INIT[579*9 +: 8], INIT[578*9 +: 8], INIT[577*9 +: 8], INIT[576*9 +: 8]}),
.INIT_13({INIT[639*9 +: 8], INIT[638*9 +: 8], INIT[637*9 +: 8], INIT[636*9 +: 8], 
          INIT[635*9 +: 8], INIT[634*9 +: 8], INIT[633*9 +: 8], INIT[632*9 +: 8], 
          INIT[631*9 +: 8], INIT[630*9 +: 8], INIT[629*9 +: 8], INIT[628*9 +: 8], 
          INIT[627*9 +: 8], INIT[626*9 +: 8], INIT[625*9 +: 8], INIT[624*9 +: 8], 
          INIT[623*9 +: 8], INIT[622*9 +: 8], INIT[621*9 +: 8], INIT[620*9 +: 8], 
          INIT[619*9 +: 8], INIT[618*9 +: 8], INIT[617*9 +: 8], INIT[616*9 +: 8], 
          INIT[615*9 +: 8], INIT[614*9 +: 8], INIT[613*9 +: 8], INIT[612*9 +: 8], 
          INIT[611*9 +: 8], INIT[610*9 +: 8], INIT[609*9 +: 8], INIT[608*9 +: 8]}),
.INIT_14({INIT[671*9 +: 8], INIT[670*9 +: 8], INIT[669*9 +: 8], INIT[668*9 +: 8], 
          INIT[667*9 +: 8], INIT[666*9 +: 8], INIT[665*9 +: 8], INIT[664*9 +: 8], 
          INIT[663*9 +: 8], INIT[662*9 +: 8], INIT[661*9 +: 8], INIT[660*9 +: 8], 
          INIT[659*9 +: 8], INIT[658*9 +: 8], INIT[657*9 +: 8], INIT[656*9 +: 8], 
          INIT[655*9 +: 8], INIT[654*9 +: 8], INIT[653*9 +: 8], INIT[652*9 +: 8], 
          INIT[651*9 +: 8], INIT[650*9 +: 8], INIT[649*9 +: 8], INIT[648*9 +: 8], 
          INIT[647*9 +: 8], INIT[646*9 +: 8], INIT[645*9 +: 8], INIT[644*9 +: 8], 
          INIT[643*9 +: 8], INIT[642*9 +: 8], INIT[641*9 +: 8], INIT[640*9 +: 8]}),
.INIT_15({INIT[703*9 +: 8], INIT[702*9 +: 8], INIT[701*9 +: 8], INIT[700*9 +: 8], 
          INIT[699*9 +: 8], INIT[698*9 +: 8], INIT[697*9 +: 8], INIT[696*9 +: 8], 
          INIT[695*9 +: 8], INIT[694*9 +: 8], INIT[693*9 +: 8], INIT[692*9 +: 8], 
          INIT[691*9 +: 8], INIT[690*9 +: 8], INIT[689*9 +: 8], INIT[688*9 +: 8], 
          INIT[687*9 +: 8], INIT[686*9 +: 8], INIT[685*9 +: 8], INIT[684*9 +: 8], 
          INIT[683*9 +: 8], INIT[682*9 +: 8], INIT[681*9 +: 8], INIT[680*9 +: 8], 
          INIT[679*9 +: 8], INIT[678*9 +: 8], INIT[677*9 +: 8], INIT[676*9 +: 8], 
          INIT[675*9 +: 8], INIT[674*9 +: 8], INIT[673*9 +: 8], INIT[672*9 +: 8]}),
.INIT_16({INIT[735*9 +: 8], INIT[734*9 +: 8], INIT[733*9 +: 8], INIT[732*9 +: 8], 
          INIT[731*9 +: 8], INIT[730*9 +: 8], INIT[729*9 +: 8], INIT[728*9 +: 8], 
          INIT[727*9 +: 8], INIT[726*9 +: 8], INIT[725*9 +: 8], INIT[724*9 +: 8], 
          INIT[723*9 +: 8], INIT[722*9 +: 8], INIT[721*9 +: 8], INIT[720*9 +: 8], 
          INIT[719*9 +: 8], INIT[718*9 +: 8], INIT[717*9 +: 8], INIT[716*9 +: 8], 
          INIT[715*9 +: 8], INIT[714*9 +: 8], INIT[713*9 +: 8], INIT[712*9 +: 8], 
          INIT[711*9 +: 8], INIT[710*9 +: 8], INIT[709*9 +: 8], INIT[708*9 +: 8], 
          INIT[707*9 +: 8], INIT[706*9 +: 8], INIT[705*9 +: 8], INIT[704*9 +: 8]}),
.INIT_17({INIT[767*9 +: 8], INIT[766*9 +: 8], INIT[765*9 +: 8], INIT[764*9 +: 8], 
          INIT[763*9 +: 8], INIT[762*9 +: 8], INIT[761*9 +: 8], INIT[760*9 +: 8], 
          INIT[759*9 +: 8], INIT[758*9 +: 8], INIT[757*9 +: 8], INIT[756*9 +: 8], 
          INIT[755*9 +: 8], INIT[754*9 +: 8], INIT[753*9 +: 8], INIT[752*9 +: 8], 
          INIT[751*9 +: 8], INIT[750*9 +: 8], INIT[749*9 +: 8], INIT[748*9 +: 8], 
          INIT[747*9 +: 8], INIT[746*9 +: 8], INIT[745*9 +: 8], INIT[744*9 +: 8], 
          INIT[743*9 +: 8], INIT[742*9 +: 8], INIT[741*9 +: 8], INIT[740*9 +: 8], 
          INIT[739*9 +: 8], INIT[738*9 +: 8], INIT[737*9 +: 8], INIT[736*9 +: 8]}),
.INIT_18({INIT[799*9 +: 8], INIT[798*9 +: 8], INIT[797*9 +: 8], INIT[796*9 +: 8], 
          INIT[795*9 +: 8], INIT[794*9 +: 8], INIT[793*9 +: 8], INIT[792*9 +: 8], 
          INIT[791*9 +: 8], INIT[790*9 +: 8], INIT[789*9 +: 8], INIT[788*9 +: 8], 
          INIT[787*9 +: 8], INIT[786*9 +: 8], INIT[785*9 +: 8], INIT[784*9 +: 8], 
          INIT[783*9 +: 8], INIT[782*9 +: 8], INIT[781*9 +: 8], INIT[780*9 +: 8], 
          INIT[779*9 +: 8], INIT[778*9 +: 8], INIT[777*9 +: 8], INIT[776*9 +: 8], 
          INIT[775*9 +: 8], INIT[774*9 +: 8], INIT[773*9 +: 8], INIT[772*9 +: 8], 
          INIT[771*9 +: 8], INIT[770*9 +: 8], INIT[769*9 +: 8], INIT[768*9 +: 8]}),
.INIT_19({INIT[831*9 +: 8], INIT[830*9 +: 8], INIT[829*9 +: 8], INIT[828*9 +: 8], 
          INIT[827*9 +: 8], INIT[826*9 +: 8], INIT[825*9 +: 8], INIT[824*9 +: 8], 
          INIT[823*9 +: 8], INIT[822*9 +: 8], INIT[821*9 +: 8], INIT[820*9 +: 8], 
          INIT[819*9 +: 8], INIT[818*9 +: 8], INIT[817*9 +: 8], INIT[816*9 +: 8], 
          INIT[815*9 +: 8], INIT[814*9 +: 8], INIT[813*9 +: 8], INIT[812*9 +: 8], 
          INIT[811*9 +: 8], INIT[810*9 +: 8], INIT[809*9 +: 8], INIT[808*9 +: 8], 
          INIT[807*9 +: 8], INIT[806*9 +: 8], INIT[805*9 +: 8], INIT[804*9 +: 8], 
          INIT[803*9 +: 8], INIT[802*9 +: 8], INIT[801*9 +: 8], INIT[800*9 +: 8]}),
.INIT_1A({INIT[863*9 +: 8], INIT[862*9 +: 8], INIT[861*9 +: 8], INIT[860*9 +: 8], 
          INIT[859*9 +: 8], INIT[858*9 +: 8], INIT[857*9 +: 8], INIT[856*9 +: 8], 
          INIT[855*9 +: 8], INIT[854*9 +: 8], INIT[853*9 +: 8], INIT[852*9 +: 8], 
          INIT[851*9 +: 8], INIT[850*9 +: 8], INIT[849*9 +: 8], INIT[848*9 +: 8], 
          INIT[847*9 +: 8], INIT[846*9 +: 8], INIT[845*9 +: 8], INIT[844*9 +: 8], 
          INIT[843*9 +: 8], INIT[842*9 +: 8], INIT[841*9 +: 8], INIT[840*9 +: 8], 
          INIT[839*9 +: 8], INIT[838*9 +: 8], INIT[837*9 +: 8], INIT[836*9 +: 8], 
          INIT[835*9 +: 8], INIT[834*9 +: 8], INIT[833*9 +: 8], INIT[832*9 +: 8]}),
.INIT_1B({INIT[895*9 +: 8], INIT[894*9 +: 8], INIT[893*9 +: 8], INIT[892*9 +: 8], 
          INIT[891*9 +: 8], INIT[890*9 +: 8], INIT[889*9 +: 8], INIT[888*9 +: 8], 
          INIT[887*9 +: 8], INIT[886*9 +: 8], INIT[885*9 +: 8], INIT[884*9 +: 8], 
          INIT[883*9 +: 8], INIT[882*9 +: 8], INIT[881*9 +: 8], INIT[880*9 +: 8], 
          INIT[879*9 +: 8], INIT[878*9 +: 8], INIT[877*9 +: 8], INIT[876*9 +: 8], 
          INIT[875*9 +: 8], INIT[874*9 +: 8], INIT[873*9 +: 8], INIT[872*9 +: 8], 
          INIT[871*9 +: 8], INIT[870*9 +: 8], INIT[869*9 +: 8], INIT[868*9 +: 8], 
          INIT[867*9 +: 8], INIT[866*9 +: 8], INIT[865*9 +: 8], INIT[864*9 +: 8]}),
.INIT_1C({INIT[927*9 +: 8], INIT[926*9 +: 8], INIT[925*9 +: 8], INIT[924*9 +: 8], 
          INIT[923*9 +: 8], INIT[922*9 +: 8], INIT[921*9 +: 8], INIT[920*9 +: 8], 
          INIT[919*9 +: 8], INIT[918*9 +: 8], INIT[917*9 +: 8], INIT[916*9 +: 8], 
          INIT[915*9 +: 8], INIT[914*9 +: 8], INIT[913*9 +: 8], INIT[912*9 +: 8], 
          INIT[911*9 +: 8], INIT[910*9 +: 8], INIT[909*9 +: 8], INIT[908*9 +: 8], 
          INIT[907*9 +: 8], INIT[906*9 +: 8], INIT[905*9 +: 8], INIT[904*9 +: 8], 
          INIT[903*9 +: 8], INIT[902*9 +: 8], INIT[901*9 +: 8], INIT[900*9 +: 8], 
          INIT[899*9 +: 8], INIT[898*9 +: 8], INIT[897*9 +: 8], INIT[896*9 +: 8]}),
.INIT_1D({INIT[959*9 +: 8], INIT[958*9 +: 8], INIT[957*9 +: 8], INIT[956*9 +: 8], 
          INIT[955*9 +: 8], INIT[954*9 +: 8], INIT[953*9 +: 8], INIT[952*9 +: 8], 
          INIT[951*9 +: 8], INIT[950*9 +: 8], INIT[949*9 +: 8], INIT[948*9 +: 8], 
          INIT[947*9 +: 8], INIT[946*9 +: 8], INIT[945*9 +: 8], INIT[944*9 +: 8], 
          INIT[943*9 +: 8], INIT[942*9 +: 8], INIT[941*9 +: 8], INIT[940*9 +: 8], 
          INIT[939*9 +: 8], INIT[938*9 +: 8], INIT[937*9 +: 8], INIT[936*9 +: 8], 
          INIT[935*9 +: 8], INIT[934*9 +: 8], INIT[933*9 +: 8], INIT[932*9 +: 8], 
          INIT[931*9 +: 8], INIT[930*9 +: 8], INIT[929*9 +: 8], INIT[928*9 +: 8]}),
.INIT_1E({INIT[991*9 +: 8], INIT[990*9 +: 8], INIT[989*9 +: 8], INIT[988*9 +: 8], 
          INIT[987*9 +: 8], INIT[986*9 +: 8], INIT[985*9 +: 8], INIT[984*9 +: 8], 
          INIT[983*9 +: 8], INIT[982*9 +: 8], INIT[981*9 +: 8], INIT[980*9 +: 8], 
          INIT[979*9 +: 8], INIT[978*9 +: 8], INIT[977*9 +: 8], INIT[976*9 +: 8], 
          INIT[975*9 +: 8], INIT[974*9 +: 8], INIT[973*9 +: 8], INIT[972*9 +: 8], 
          INIT[971*9 +: 8], INIT[970*9 +: 8], INIT[969*9 +: 8], INIT[968*9 +: 8], 
          INIT[967*9 +: 8], INIT[966*9 +: 8], INIT[965*9 +: 8], INIT[964*9 +: 8], 
          INIT[963*9 +: 8], INIT[962*9 +: 8], INIT[961*9 +: 8], INIT[960*9 +: 8]}),
.INIT_1F({INIT[1023*9 +: 8], INIT[1022*9 +: 8], INIT[1021*9 +: 8], INIT[1020*9 +: 8], 
          INIT[1019*9 +: 8], INIT[1018*9 +: 8], INIT[1017*9 +: 8], INIT[1016*9 +: 8], 
          INIT[1015*9 +: 8], INIT[1014*9 +: 8], INIT[1013*9 +: 8], INIT[1012*9 +: 8], 
          INIT[1011*9 +: 8], INIT[1010*9 +: 8], INIT[1009*9 +: 8], INIT[1008*9 +: 8], 
          INIT[1007*9 +: 8], INIT[1006*9 +: 8], INIT[1005*9 +: 8], INIT[1004*9 +: 8], 
          INIT[1003*9 +: 8], INIT[1002*9 +: 8], INIT[1001*9 +: 8], INIT[1000*9 +: 8], 
          INIT[999*9 +: 8], INIT[998*9 +: 8], INIT[997*9 +: 8], INIT[996*9 +: 8], 
          INIT[995*9 +: 8], INIT[994*9 +: 8], INIT[993*9 +: 8], INIT[992*9 +: 8]}),
.INIT_20({INIT[1055*9 +: 8], INIT[1054*9 +: 8], INIT[1053*9 +: 8], INIT[1052*9 +: 8], 
          INIT[1051*9 +: 8], INIT[1050*9 +: 8], INIT[1049*9 +: 8], INIT[1048*9 +: 8], 
          INIT[1047*9 +: 8], INIT[1046*9 +: 8], INIT[1045*9 +: 8], INIT[1044*9 +: 8], 
          INIT[1043*9 +: 8], INIT[1042*9 +: 8], INIT[1041*9 +: 8], INIT[1040*9 +: 8], 
          INIT[1039*9 +: 8], INIT[1038*9 +: 8], INIT[1037*9 +: 8], INIT[1036*9 +: 8], 
          INIT[1035*9 +: 8], INIT[1034*9 +: 8], INIT[1033*9 +: 8], INIT[1032*9 +: 8], 
          INIT[1031*9 +: 8], INIT[1030*9 +: 8], INIT[1029*9 +: 8], INIT[1028*9 +: 8], 
          INIT[1027*9 +: 8], INIT[1026*9 +: 8], INIT[1025*9 +: 8], INIT[1024*9 +: 8]}),
.INIT_21({INIT[1087*9 +: 8], INIT[1086*9 +: 8], INIT[1085*9 +: 8], INIT[1084*9 +: 8], 
          INIT[1083*9 +: 8], INIT[1082*9 +: 8], INIT[1081*9 +: 8], INIT[1080*9 +: 8], 
          INIT[1079*9 +: 8], INIT[1078*9 +: 8], INIT[1077*9 +: 8], INIT[1076*9 +: 8], 
          INIT[1075*9 +: 8], INIT[1074*9 +: 8], INIT[1073*9 +: 8], INIT[1072*9 +: 8], 
          INIT[1071*9 +: 8], INIT[1070*9 +: 8], INIT[1069*9 +: 8], INIT[1068*9 +: 8], 
          INIT[1067*9 +: 8], INIT[1066*9 +: 8], INIT[1065*9 +: 8], INIT[1064*9 +: 8], 
          INIT[1063*9 +: 8], INIT[1062*9 +: 8], INIT[1061*9 +: 8], INIT[1060*9 +: 8], 
          INIT[1059*9 +: 8], INIT[1058*9 +: 8], INIT[1057*9 +: 8], INIT[1056*9 +: 8]}),
.INIT_22({INIT[1119*9 +: 8], INIT[1118*9 +: 8], INIT[1117*9 +: 8], INIT[1116*9 +: 8], 
          INIT[1115*9 +: 8], INIT[1114*9 +: 8], INIT[1113*9 +: 8], INIT[1112*9 +: 8], 
          INIT[1111*9 +: 8], INIT[1110*9 +: 8], INIT[1109*9 +: 8], INIT[1108*9 +: 8], 
          INIT[1107*9 +: 8], INIT[1106*9 +: 8], INIT[1105*9 +: 8], INIT[1104*9 +: 8], 
          INIT[1103*9 +: 8], INIT[1102*9 +: 8], INIT[1101*9 +: 8], INIT[1100*9 +: 8], 
          INIT[1099*9 +: 8], INIT[1098*9 +: 8], INIT[1097*9 +: 8], INIT[1096*9 +: 8], 
          INIT[1095*9 +: 8], INIT[1094*9 +: 8], INIT[1093*9 +: 8], INIT[1092*9 +: 8], 
          INIT[1091*9 +: 8], INIT[1090*9 +: 8], INIT[1089*9 +: 8], INIT[1088*9 +: 8]}),
.INIT_23({INIT[1151*9 +: 8], INIT[1150*9 +: 8], INIT[1149*9 +: 8], INIT[1148*9 +: 8], 
          INIT[1147*9 +: 8], INIT[1146*9 +: 8], INIT[1145*9 +: 8], INIT[1144*9 +: 8], 
          INIT[1143*9 +: 8], INIT[1142*9 +: 8], INIT[1141*9 +: 8], INIT[1140*9 +: 8], 
          INIT[1139*9 +: 8], INIT[1138*9 +: 8], INIT[1137*9 +: 8], INIT[1136*9 +: 8], 
          INIT[1135*9 +: 8], INIT[1134*9 +: 8], INIT[1133*9 +: 8], INIT[1132*9 +: 8], 
          INIT[1131*9 +: 8], INIT[1130*9 +: 8], INIT[1129*9 +: 8], INIT[1128*9 +: 8], 
          INIT[1127*9 +: 8], INIT[1126*9 +: 8], INIT[1125*9 +: 8], INIT[1124*9 +: 8], 
          INIT[1123*9 +: 8], INIT[1122*9 +: 8], INIT[1121*9 +: 8], INIT[1120*9 +: 8]}),
.INIT_24({INIT[1183*9 +: 8], INIT[1182*9 +: 8], INIT[1181*9 +: 8], INIT[1180*9 +: 8], 
          INIT[1179*9 +: 8], INIT[1178*9 +: 8], INIT[1177*9 +: 8], INIT[1176*9 +: 8], 
          INIT[1175*9 +: 8], INIT[1174*9 +: 8], INIT[1173*9 +: 8], INIT[1172*9 +: 8], 
          INIT[1171*9 +: 8], INIT[1170*9 +: 8], INIT[1169*9 +: 8], INIT[1168*9 +: 8], 
          INIT[1167*9 +: 8], INIT[1166*9 +: 8], INIT[1165*9 +: 8], INIT[1164*9 +: 8], 
          INIT[1163*9 +: 8], INIT[1162*9 +: 8], INIT[1161*9 +: 8], INIT[1160*9 +: 8], 
          INIT[1159*9 +: 8], INIT[1158*9 +: 8], INIT[1157*9 +: 8], INIT[1156*9 +: 8], 
          INIT[1155*9 +: 8], INIT[1154*9 +: 8], INIT[1153*9 +: 8], INIT[1152*9 +: 8]}),
.INIT_25({INIT[1215*9 +: 8], INIT[1214*9 +: 8], INIT[1213*9 +: 8], INIT[1212*9 +: 8], 
          INIT[1211*9 +: 8], INIT[1210*9 +: 8], INIT[1209*9 +: 8], INIT[1208*9 +: 8], 
          INIT[1207*9 +: 8], INIT[1206*9 +: 8], INIT[1205*9 +: 8], INIT[1204*9 +: 8], 
          INIT[1203*9 +: 8], INIT[1202*9 +: 8], INIT[1201*9 +: 8], INIT[1200*9 +: 8], 
          INIT[1199*9 +: 8], INIT[1198*9 +: 8], INIT[1197*9 +: 8], INIT[1196*9 +: 8], 
          INIT[1195*9 +: 8], INIT[1194*9 +: 8], INIT[1193*9 +: 8], INIT[1192*9 +: 8], 
          INIT[1191*9 +: 8], INIT[1190*9 +: 8], INIT[1189*9 +: 8], INIT[1188*9 +: 8], 
          INIT[1187*9 +: 8], INIT[1186*9 +: 8], INIT[1185*9 +: 8], INIT[1184*9 +: 8]}),
.INIT_26({INIT[1247*9 +: 8], INIT[1246*9 +: 8], INIT[1245*9 +: 8], INIT[1244*9 +: 8], 
          INIT[1243*9 +: 8], INIT[1242*9 +: 8], INIT[1241*9 +: 8], INIT[1240*9 +: 8], 
          INIT[1239*9 +: 8], INIT[1238*9 +: 8], INIT[1237*9 +: 8], INIT[1236*9 +: 8], 
          INIT[1235*9 +: 8], INIT[1234*9 +: 8], INIT[1233*9 +: 8], INIT[1232*9 +: 8], 
          INIT[1231*9 +: 8], INIT[1230*9 +: 8], INIT[1229*9 +: 8], INIT[1228*9 +: 8], 
          INIT[1227*9 +: 8], INIT[1226*9 +: 8], INIT[1225*9 +: 8], INIT[1224*9 +: 8], 
          INIT[1223*9 +: 8], INIT[1222*9 +: 8], INIT[1221*9 +: 8], INIT[1220*9 +: 8], 
          INIT[1219*9 +: 8], INIT[1218*9 +: 8], INIT[1217*9 +: 8], INIT[1216*9 +: 8]}),
.INIT_27({INIT[1279*9 +: 8], INIT[1278*9 +: 8], INIT[1277*9 +: 8], INIT[1276*9 +: 8], 
          INIT[1275*9 +: 8], INIT[1274*9 +: 8], INIT[1273*9 +: 8], INIT[1272*9 +: 8], 
          INIT[1271*9 +: 8], INIT[1270*9 +: 8], INIT[1269*9 +: 8], INIT[1268*9 +: 8], 
          INIT[1267*9 +: 8], INIT[1266*9 +: 8], INIT[1265*9 +: 8], INIT[1264*9 +: 8], 
          INIT[1263*9 +: 8], INIT[1262*9 +: 8], INIT[1261*9 +: 8], INIT[1260*9 +: 8], 
          INIT[1259*9 +: 8], INIT[1258*9 +: 8], INIT[1257*9 +: 8], INIT[1256*9 +: 8], 
          INIT[1255*9 +: 8], INIT[1254*9 +: 8], INIT[1253*9 +: 8], INIT[1252*9 +: 8], 
          INIT[1251*9 +: 8], INIT[1250*9 +: 8], INIT[1249*9 +: 8], INIT[1248*9 +: 8]}),
.INIT_28({INIT[1311*9 +: 8], INIT[1310*9 +: 8], INIT[1309*9 +: 8], INIT[1308*9 +: 8], 
          INIT[1307*9 +: 8], INIT[1306*9 +: 8], INIT[1305*9 +: 8], INIT[1304*9 +: 8], 
          INIT[1303*9 +: 8], INIT[1302*9 +: 8], INIT[1301*9 +: 8], INIT[1300*9 +: 8], 
          INIT[1299*9 +: 8], INIT[1298*9 +: 8], INIT[1297*9 +: 8], INIT[1296*9 +: 8], 
          INIT[1295*9 +: 8], INIT[1294*9 +: 8], INIT[1293*9 +: 8], INIT[1292*9 +: 8], 
          INIT[1291*9 +: 8], INIT[1290*9 +: 8], INIT[1289*9 +: 8], INIT[1288*9 +: 8], 
          INIT[1287*9 +: 8], INIT[1286*9 +: 8], INIT[1285*9 +: 8], INIT[1284*9 +: 8], 
          INIT[1283*9 +: 8], INIT[1282*9 +: 8], INIT[1281*9 +: 8], INIT[1280*9 +: 8]}),
.INIT_29({INIT[1343*9 +: 8], INIT[1342*9 +: 8], INIT[1341*9 +: 8], INIT[1340*9 +: 8], 
          INIT[1339*9 +: 8], INIT[1338*9 +: 8], INIT[1337*9 +: 8], INIT[1336*9 +: 8], 
          INIT[1335*9 +: 8], INIT[1334*9 +: 8], INIT[1333*9 +: 8], INIT[1332*9 +: 8], 
          INIT[1331*9 +: 8], INIT[1330*9 +: 8], INIT[1329*9 +: 8], INIT[1328*9 +: 8], 
          INIT[1327*9 +: 8], INIT[1326*9 +: 8], INIT[1325*9 +: 8], INIT[1324*9 +: 8], 
          INIT[1323*9 +: 8], INIT[1322*9 +: 8], INIT[1321*9 +: 8], INIT[1320*9 +: 8], 
          INIT[1319*9 +: 8], INIT[1318*9 +: 8], INIT[1317*9 +: 8], INIT[1316*9 +: 8], 
          INIT[1315*9 +: 8], INIT[1314*9 +: 8], INIT[1313*9 +: 8], INIT[1312*9 +: 8]}),
.INIT_2A({INIT[1375*9 +: 8], INIT[1374*9 +: 8], INIT[1373*9 +: 8], INIT[1372*9 +: 8], 
          INIT[1371*9 +: 8], INIT[1370*9 +: 8], INIT[1369*9 +: 8], INIT[1368*9 +: 8], 
          INIT[1367*9 +: 8], INIT[1366*9 +: 8], INIT[1365*9 +: 8], INIT[1364*9 +: 8], 
          INIT[1363*9 +: 8], INIT[1362*9 +: 8], INIT[1361*9 +: 8], INIT[1360*9 +: 8], 
          INIT[1359*9 +: 8], INIT[1358*9 +: 8], INIT[1357*9 +: 8], INIT[1356*9 +: 8], 
          INIT[1355*9 +: 8], INIT[1354*9 +: 8], INIT[1353*9 +: 8], INIT[1352*9 +: 8], 
          INIT[1351*9 +: 8], INIT[1350*9 +: 8], INIT[1349*9 +: 8], INIT[1348*9 +: 8], 
          INIT[1347*9 +: 8], INIT[1346*9 +: 8], INIT[1345*9 +: 8], INIT[1344*9 +: 8]}),
.INIT_2B({INIT[1407*9 +: 8], INIT[1406*9 +: 8], INIT[1405*9 +: 8], INIT[1404*9 +: 8], 
          INIT[1403*9 +: 8], INIT[1402*9 +: 8], INIT[1401*9 +: 8], INIT[1400*9 +: 8], 
          INIT[1399*9 +: 8], INIT[1398*9 +: 8], INIT[1397*9 +: 8], INIT[1396*9 +: 8], 
          INIT[1395*9 +: 8], INIT[1394*9 +: 8], INIT[1393*9 +: 8], INIT[1392*9 +: 8], 
          INIT[1391*9 +: 8], INIT[1390*9 +: 8], INIT[1389*9 +: 8], INIT[1388*9 +: 8], 
          INIT[1387*9 +: 8], INIT[1386*9 +: 8], INIT[1385*9 +: 8], INIT[1384*9 +: 8], 
          INIT[1383*9 +: 8], INIT[1382*9 +: 8], INIT[1381*9 +: 8], INIT[1380*9 +: 8], 
          INIT[1379*9 +: 8], INIT[1378*9 +: 8], INIT[1377*9 +: 8], INIT[1376*9 +: 8]}),
.INIT_2C({INIT[1439*9 +: 8], INIT[1438*9 +: 8], INIT[1437*9 +: 8], INIT[1436*9 +: 8], 
          INIT[1435*9 +: 8], INIT[1434*9 +: 8], INIT[1433*9 +: 8], INIT[1432*9 +: 8], 
          INIT[1431*9 +: 8], INIT[1430*9 +: 8], INIT[1429*9 +: 8], INIT[1428*9 +: 8], 
          INIT[1427*9 +: 8], INIT[1426*9 +: 8], INIT[1425*9 +: 8], INIT[1424*9 +: 8], 
          INIT[1423*9 +: 8], INIT[1422*9 +: 8], INIT[1421*9 +: 8], INIT[1420*9 +: 8], 
          INIT[1419*9 +: 8], INIT[1418*9 +: 8], INIT[1417*9 +: 8], INIT[1416*9 +: 8], 
          INIT[1415*9 +: 8], INIT[1414*9 +: 8], INIT[1413*9 +: 8], INIT[1412*9 +: 8], 
          INIT[1411*9 +: 8], INIT[1410*9 +: 8], INIT[1409*9 +: 8], INIT[1408*9 +: 8]}),
.INIT_2D({INIT[1471*9 +: 8], INIT[1470*9 +: 8], INIT[1469*9 +: 8], INIT[1468*9 +: 8], 
          INIT[1467*9 +: 8], INIT[1466*9 +: 8], INIT[1465*9 +: 8], INIT[1464*9 +: 8], 
          INIT[1463*9 +: 8], INIT[1462*9 +: 8], INIT[1461*9 +: 8], INIT[1460*9 +: 8], 
          INIT[1459*9 +: 8], INIT[1458*9 +: 8], INIT[1457*9 +: 8], INIT[1456*9 +: 8], 
          INIT[1455*9 +: 8], INIT[1454*9 +: 8], INIT[1453*9 +: 8], INIT[1452*9 +: 8], 
          INIT[1451*9 +: 8], INIT[1450*9 +: 8], INIT[1449*9 +: 8], INIT[1448*9 +: 8], 
          INIT[1447*9 +: 8], INIT[1446*9 +: 8], INIT[1445*9 +: 8], INIT[1444*9 +: 8], 
          INIT[1443*9 +: 8], INIT[1442*9 +: 8], INIT[1441*9 +: 8], INIT[1440*9 +: 8]}),
.INIT_2E({INIT[1503*9 +: 8], INIT[1502*9 +: 8], INIT[1501*9 +: 8], INIT[1500*9 +: 8], 
          INIT[1499*9 +: 8], INIT[1498*9 +: 8], INIT[1497*9 +: 8], INIT[1496*9 +: 8], 
          INIT[1495*9 +: 8], INIT[1494*9 +: 8], INIT[1493*9 +: 8], INIT[1492*9 +: 8], 
          INIT[1491*9 +: 8], INIT[1490*9 +: 8], INIT[1489*9 +: 8], INIT[1488*9 +: 8], 
          INIT[1487*9 +: 8], INIT[1486*9 +: 8], INIT[1485*9 +: 8], INIT[1484*9 +: 8], 
          INIT[1483*9 +: 8], INIT[1482*9 +: 8], INIT[1481*9 +: 8], INIT[1480*9 +: 8], 
          INIT[1479*9 +: 8], INIT[1478*9 +: 8], INIT[1477*9 +: 8], INIT[1476*9 +: 8], 
          INIT[1475*9 +: 8], INIT[1474*9 +: 8], INIT[1473*9 +: 8], INIT[1472*9 +: 8]}),
.INIT_2F({INIT[1535*9 +: 8], INIT[1534*9 +: 8], INIT[1533*9 +: 8], INIT[1532*9 +: 8], 
          INIT[1531*9 +: 8], INIT[1530*9 +: 8], INIT[1529*9 +: 8], INIT[1528*9 +: 8], 
          INIT[1527*9 +: 8], INIT[1526*9 +: 8], INIT[1525*9 +: 8], INIT[1524*9 +: 8], 
          INIT[1523*9 +: 8], INIT[1522*9 +: 8], INIT[1521*9 +: 8], INIT[1520*9 +: 8], 
          INIT[1519*9 +: 8], INIT[1518*9 +: 8], INIT[1517*9 +: 8], INIT[1516*9 +: 8], 
          INIT[1515*9 +: 8], INIT[1514*9 +: 8], INIT[1513*9 +: 8], INIT[1512*9 +: 8], 
          INIT[1511*9 +: 8], INIT[1510*9 +: 8], INIT[1509*9 +: 8], INIT[1508*9 +: 8], 
          INIT[1507*9 +: 8], INIT[1506*9 +: 8], INIT[1505*9 +: 8], INIT[1504*9 +: 8]}),
.INIT_30({INIT[1567*9 +: 8], INIT[1566*9 +: 8], INIT[1565*9 +: 8], INIT[1564*9 +: 8], 
          INIT[1563*9 +: 8], INIT[1562*9 +: 8], INIT[1561*9 +: 8], INIT[1560*9 +: 8], 
          INIT[1559*9 +: 8], INIT[1558*9 +: 8], INIT[1557*9 +: 8], INIT[1556*9 +: 8], 
          INIT[1555*9 +: 8], INIT[1554*9 +: 8], INIT[1553*9 +: 8], INIT[1552*9 +: 8], 
          INIT[1551*9 +: 8], INIT[1550*9 +: 8], INIT[1549*9 +: 8], INIT[1548*9 +: 8], 
          INIT[1547*9 +: 8], INIT[1546*9 +: 8], INIT[1545*9 +: 8], INIT[1544*9 +: 8], 
          INIT[1543*9 +: 8], INIT[1542*9 +: 8], INIT[1541*9 +: 8], INIT[1540*9 +: 8], 
          INIT[1539*9 +: 8], INIT[1538*9 +: 8], INIT[1537*9 +: 8], INIT[1536*9 +: 8]}),
.INIT_31({INIT[1599*9 +: 8], INIT[1598*9 +: 8], INIT[1597*9 +: 8], INIT[1596*9 +: 8], 
          INIT[1595*9 +: 8], INIT[1594*9 +: 8], INIT[1593*9 +: 8], INIT[1592*9 +: 8], 
          INIT[1591*9 +: 8], INIT[1590*9 +: 8], INIT[1589*9 +: 8], INIT[1588*9 +: 8], 
          INIT[1587*9 +: 8], INIT[1586*9 +: 8], INIT[1585*9 +: 8], INIT[1584*9 +: 8], 
          INIT[1583*9 +: 8], INIT[1582*9 +: 8], INIT[1581*9 +: 8], INIT[1580*9 +: 8], 
          INIT[1579*9 +: 8], INIT[1578*9 +: 8], INIT[1577*9 +: 8], INIT[1576*9 +: 8], 
          INIT[1575*9 +: 8], INIT[1574*9 +: 8], INIT[1573*9 +: 8], INIT[1572*9 +: 8], 
          INIT[1571*9 +: 8], INIT[1570*9 +: 8], INIT[1569*9 +: 8], INIT[1568*9 +: 8]}),
.INIT_32({INIT[1631*9 +: 8], INIT[1630*9 +: 8], INIT[1629*9 +: 8], INIT[1628*9 +: 8], 
          INIT[1627*9 +: 8], INIT[1626*9 +: 8], INIT[1625*9 +: 8], INIT[1624*9 +: 8], 
          INIT[1623*9 +: 8], INIT[1622*9 +: 8], INIT[1621*9 +: 8], INIT[1620*9 +: 8], 
          INIT[1619*9 +: 8], INIT[1618*9 +: 8], INIT[1617*9 +: 8], INIT[1616*9 +: 8], 
          INIT[1615*9 +: 8], INIT[1614*9 +: 8], INIT[1613*9 +: 8], INIT[1612*9 +: 8], 
          INIT[1611*9 +: 8], INIT[1610*9 +: 8], INIT[1609*9 +: 8], INIT[1608*9 +: 8], 
          INIT[1607*9 +: 8], INIT[1606*9 +: 8], INIT[1605*9 +: 8], INIT[1604*9 +: 8], 
          INIT[1603*9 +: 8], INIT[1602*9 +: 8], INIT[1601*9 +: 8], INIT[1600*9 +: 8]}),
.INIT_33({INIT[1663*9 +: 8], INIT[1662*9 +: 8], INIT[1661*9 +: 8], INIT[1660*9 +: 8], 
          INIT[1659*9 +: 8], INIT[1658*9 +: 8], INIT[1657*9 +: 8], INIT[1656*9 +: 8], 
          INIT[1655*9 +: 8], INIT[1654*9 +: 8], INIT[1653*9 +: 8], INIT[1652*9 +: 8], 
          INIT[1651*9 +: 8], INIT[1650*9 +: 8], INIT[1649*9 +: 8], INIT[1648*9 +: 8], 
          INIT[1647*9 +: 8], INIT[1646*9 +: 8], INIT[1645*9 +: 8], INIT[1644*9 +: 8], 
          INIT[1643*9 +: 8], INIT[1642*9 +: 8], INIT[1641*9 +: 8], INIT[1640*9 +: 8], 
          INIT[1639*9 +: 8], INIT[1638*9 +: 8], INIT[1637*9 +: 8], INIT[1636*9 +: 8], 
          INIT[1635*9 +: 8], INIT[1634*9 +: 8], INIT[1633*9 +: 8], INIT[1632*9 +: 8]}),
.INIT_34({INIT[1695*9 +: 8], INIT[1694*9 +: 8], INIT[1693*9 +: 8], INIT[1692*9 +: 8], 
          INIT[1691*9 +: 8], INIT[1690*9 +: 8], INIT[1689*9 +: 8], INIT[1688*9 +: 8], 
          INIT[1687*9 +: 8], INIT[1686*9 +: 8], INIT[1685*9 +: 8], INIT[1684*9 +: 8], 
          INIT[1683*9 +: 8], INIT[1682*9 +: 8], INIT[1681*9 +: 8], INIT[1680*9 +: 8], 
          INIT[1679*9 +: 8], INIT[1678*9 +: 8], INIT[1677*9 +: 8], INIT[1676*9 +: 8], 
          INIT[1675*9 +: 8], INIT[1674*9 +: 8], INIT[1673*9 +: 8], INIT[1672*9 +: 8], 
          INIT[1671*9 +: 8], INIT[1670*9 +: 8], INIT[1669*9 +: 8], INIT[1668*9 +: 8], 
          INIT[1667*9 +: 8], INIT[1666*9 +: 8], INIT[1665*9 +: 8], INIT[1664*9 +: 8]}),
.INIT_35({INIT[1727*9 +: 8], INIT[1726*9 +: 8], INIT[1725*9 +: 8], INIT[1724*9 +: 8], 
          INIT[1723*9 +: 8], INIT[1722*9 +: 8], INIT[1721*9 +: 8], INIT[1720*9 +: 8], 
          INIT[1719*9 +: 8], INIT[1718*9 +: 8], INIT[1717*9 +: 8], INIT[1716*9 +: 8], 
          INIT[1715*9 +: 8], INIT[1714*9 +: 8], INIT[1713*9 +: 8], INIT[1712*9 +: 8], 
          INIT[1711*9 +: 8], INIT[1710*9 +: 8], INIT[1709*9 +: 8], INIT[1708*9 +: 8], 
          INIT[1707*9 +: 8], INIT[1706*9 +: 8], INIT[1705*9 +: 8], INIT[1704*9 +: 8], 
          INIT[1703*9 +: 8], INIT[1702*9 +: 8], INIT[1701*9 +: 8], INIT[1700*9 +: 8], 
          INIT[1699*9 +: 8], INIT[1698*9 +: 8], INIT[1697*9 +: 8], INIT[1696*9 +: 8]}),
.INIT_36({INIT[1759*9 +: 8], INIT[1758*9 +: 8], INIT[1757*9 +: 8], INIT[1756*9 +: 8], 
          INIT[1755*9 +: 8], INIT[1754*9 +: 8], INIT[1753*9 +: 8], INIT[1752*9 +: 8], 
          INIT[1751*9 +: 8], INIT[1750*9 +: 8], INIT[1749*9 +: 8], INIT[1748*9 +: 8], 
          INIT[1747*9 +: 8], INIT[1746*9 +: 8], INIT[1745*9 +: 8], INIT[1744*9 +: 8], 
          INIT[1743*9 +: 8], INIT[1742*9 +: 8], INIT[1741*9 +: 8], INIT[1740*9 +: 8], 
          INIT[1739*9 +: 8], INIT[1738*9 +: 8], INIT[1737*9 +: 8], INIT[1736*9 +: 8], 
          INIT[1735*9 +: 8], INIT[1734*9 +: 8], INIT[1733*9 +: 8], INIT[1732*9 +: 8], 
          INIT[1731*9 +: 8], INIT[1730*9 +: 8], INIT[1729*9 +: 8], INIT[1728*9 +: 8]}),
.INIT_37({INIT[1791*9 +: 8], INIT[1790*9 +: 8], INIT[1789*9 +: 8], INIT[1788*9 +: 8], 
          INIT[1787*9 +: 8], INIT[1786*9 +: 8], INIT[1785*9 +: 8], INIT[1784*9 +: 8], 
          INIT[1783*9 +: 8], INIT[1782*9 +: 8], INIT[1781*9 +: 8], INIT[1780*9 +: 8], 
          INIT[1779*9 +: 8], INIT[1778*9 +: 8], INIT[1777*9 +: 8], INIT[1776*9 +: 8], 
          INIT[1775*9 +: 8], INIT[1774*9 +: 8], INIT[1773*9 +: 8], INIT[1772*9 +: 8], 
          INIT[1771*9 +: 8], INIT[1770*9 +: 8], INIT[1769*9 +: 8], INIT[1768*9 +: 8], 
          INIT[1767*9 +: 8], INIT[1766*9 +: 8], INIT[1765*9 +: 8], INIT[1764*9 +: 8], 
          INIT[1763*9 +: 8], INIT[1762*9 +: 8], INIT[1761*9 +: 8], INIT[1760*9 +: 8]}),
.INIT_38({INIT[1823*9 +: 8], INIT[1822*9 +: 8], INIT[1821*9 +: 8], INIT[1820*9 +: 8], 
          INIT[1819*9 +: 8], INIT[1818*9 +: 8], INIT[1817*9 +: 8], INIT[1816*9 +: 8], 
          INIT[1815*9 +: 8], INIT[1814*9 +: 8], INIT[1813*9 +: 8], INIT[1812*9 +: 8], 
          INIT[1811*9 +: 8], INIT[1810*9 +: 8], INIT[1809*9 +: 8], INIT[1808*9 +: 8], 
          INIT[1807*9 +: 8], INIT[1806*9 +: 8], INIT[1805*9 +: 8], INIT[1804*9 +: 8], 
          INIT[1803*9 +: 8], INIT[1802*9 +: 8], INIT[1801*9 +: 8], INIT[1800*9 +: 8], 
          INIT[1799*9 +: 8], INIT[1798*9 +: 8], INIT[1797*9 +: 8], INIT[1796*9 +: 8], 
          INIT[1795*9 +: 8], INIT[1794*9 +: 8], INIT[1793*9 +: 8], INIT[1792*9 +: 8]}),
.INIT_39({INIT[1855*9 +: 8], INIT[1854*9 +: 8], INIT[1853*9 +: 8], INIT[1852*9 +: 8], 
          INIT[1851*9 +: 8], INIT[1850*9 +: 8], INIT[1849*9 +: 8], INIT[1848*9 +: 8], 
          INIT[1847*9 +: 8], INIT[1846*9 +: 8], INIT[1845*9 +: 8], INIT[1844*9 +: 8], 
          INIT[1843*9 +: 8], INIT[1842*9 +: 8], INIT[1841*9 +: 8], INIT[1840*9 +: 8], 
          INIT[1839*9 +: 8], INIT[1838*9 +: 8], INIT[1837*9 +: 8], INIT[1836*9 +: 8], 
          INIT[1835*9 +: 8], INIT[1834*9 +: 8], INIT[1833*9 +: 8], INIT[1832*9 +: 8], 
          INIT[1831*9 +: 8], INIT[1830*9 +: 8], INIT[1829*9 +: 8], INIT[1828*9 +: 8], 
          INIT[1827*9 +: 8], INIT[1826*9 +: 8], INIT[1825*9 +: 8], INIT[1824*9 +: 8]}),
.INIT_3A({INIT[1887*9 +: 8], INIT[1886*9 +: 8], INIT[1885*9 +: 8], INIT[1884*9 +: 8], 
          INIT[1883*9 +: 8], INIT[1882*9 +: 8], INIT[1881*9 +: 8], INIT[1880*9 +: 8], 
          INIT[1879*9 +: 8], INIT[1878*9 +: 8], INIT[1877*9 +: 8], INIT[1876*9 +: 8], 
          INIT[1875*9 +: 8], INIT[1874*9 +: 8], INIT[1873*9 +: 8], INIT[1872*9 +: 8], 
          INIT[1871*9 +: 8], INIT[1870*9 +: 8], INIT[1869*9 +: 8], INIT[1868*9 +: 8], 
          INIT[1867*9 +: 8], INIT[1866*9 +: 8], INIT[1865*9 +: 8], INIT[1864*9 +: 8], 
          INIT[1863*9 +: 8], INIT[1862*9 +: 8], INIT[1861*9 +: 8], INIT[1860*9 +: 8], 
          INIT[1859*9 +: 8], INIT[1858*9 +: 8], INIT[1857*9 +: 8], INIT[1856*9 +: 8]}),
.INIT_3B({INIT[1919*9 +: 8], INIT[1918*9 +: 8], INIT[1917*9 +: 8], INIT[1916*9 +: 8], 
          INIT[1915*9 +: 8], INIT[1914*9 +: 8], INIT[1913*9 +: 8], INIT[1912*9 +: 8], 
          INIT[1911*9 +: 8], INIT[1910*9 +: 8], INIT[1909*9 +: 8], INIT[1908*9 +: 8], 
          INIT[1907*9 +: 8], INIT[1906*9 +: 8], INIT[1905*9 +: 8], INIT[1904*9 +: 8], 
          INIT[1903*9 +: 8], INIT[1902*9 +: 8], INIT[1901*9 +: 8], INIT[1900*9 +: 8], 
          INIT[1899*9 +: 8], INIT[1898*9 +: 8], INIT[1897*9 +: 8], INIT[1896*9 +: 8], 
          INIT[1895*9 +: 8], INIT[1894*9 +: 8], INIT[1893*9 +: 8], INIT[1892*9 +: 8], 
          INIT[1891*9 +: 8], INIT[1890*9 +: 8], INIT[1889*9 +: 8], INIT[1888*9 +: 8]}),
.INIT_3C({INIT[1951*9 +: 8], INIT[1950*9 +: 8], INIT[1949*9 +: 8], INIT[1948*9 +: 8], 
          INIT[1947*9 +: 8], INIT[1946*9 +: 8], INIT[1945*9 +: 8], INIT[1944*9 +: 8], 
          INIT[1943*9 +: 8], INIT[1942*9 +: 8], INIT[1941*9 +: 8], INIT[1940*9 +: 8], 
          INIT[1939*9 +: 8], INIT[1938*9 +: 8], INIT[1937*9 +: 8], INIT[1936*9 +: 8], 
          INIT[1935*9 +: 8], INIT[1934*9 +: 8], INIT[1933*9 +: 8], INIT[1932*9 +: 8], 
          INIT[1931*9 +: 8], INIT[1930*9 +: 8], INIT[1929*9 +: 8], INIT[1928*9 +: 8], 
          INIT[1927*9 +: 8], INIT[1926*9 +: 8], INIT[1925*9 +: 8], INIT[1924*9 +: 8], 
          INIT[1923*9 +: 8], INIT[1922*9 +: 8], INIT[1921*9 +: 8], INIT[1920*9 +: 8]}),
.INIT_3D({INIT[1983*9 +: 8], INIT[1982*9 +: 8], INIT[1981*9 +: 8], INIT[1980*9 +: 8], 
          INIT[1979*9 +: 8], INIT[1978*9 +: 8], INIT[1977*9 +: 8], INIT[1976*9 +: 8], 
          INIT[1975*9 +: 8], INIT[1974*9 +: 8], INIT[1973*9 +: 8], INIT[1972*9 +: 8], 
          INIT[1971*9 +: 8], INIT[1970*9 +: 8], INIT[1969*9 +: 8], INIT[1968*9 +: 8], 
          INIT[1967*9 +: 8], INIT[1966*9 +: 8], INIT[1965*9 +: 8], INIT[1964*9 +: 8], 
          INIT[1963*9 +: 8], INIT[1962*9 +: 8], INIT[1961*9 +: 8], INIT[1960*9 +: 8], 
          INIT[1959*9 +: 8], INIT[1958*9 +: 8], INIT[1957*9 +: 8], INIT[1956*9 +: 8], 
          INIT[1955*9 +: 8], INIT[1954*9 +: 8], INIT[1953*9 +: 8], INIT[1952*9 +: 8]}),
.INIT_3E({INIT[2015*9 +: 8], INIT[2014*9 +: 8], INIT[2013*9 +: 8], INIT[2012*9 +: 8], 
          INIT[2011*9 +: 8], INIT[2010*9 +: 8], INIT[2009*9 +: 8], INIT[2008*9 +: 8], 
          INIT[2007*9 +: 8], INIT[2006*9 +: 8], INIT[2005*9 +: 8], INIT[2004*9 +: 8], 
          INIT[2003*9 +: 8], INIT[2002*9 +: 8], INIT[2001*9 +: 8], INIT[2000*9 +: 8], 
          INIT[1999*9 +: 8], INIT[1998*9 +: 8], INIT[1997*9 +: 8], INIT[1996*9 +: 8], 
          INIT[1995*9 +: 8], INIT[1994*9 +: 8], INIT[1993*9 +: 8], INIT[1992*9 +: 8], 
          INIT[1991*9 +: 8], INIT[1990*9 +: 8], INIT[1989*9 +: 8], INIT[1988*9 +: 8], 
          INIT[1987*9 +: 8], INIT[1986*9 +: 8], INIT[1985*9 +: 8], INIT[1984*9 +: 8]}),
.INIT_3F({INIT[2047*9 +: 8], INIT[2046*9 +: 8], INIT[2045*9 +: 8], INIT[2044*9 +: 8], 
          INIT[2043*9 +: 8], INIT[2042*9 +: 8], INIT[2041*9 +: 8], INIT[2040*9 +: 8], 
          INIT[2039*9 +: 8], INIT[2038*9 +: 8], INIT[2037*9 +: 8], INIT[2036*9 +: 8], 
          INIT[2035*9 +: 8], INIT[2034*9 +: 8], INIT[2033*9 +: 8], INIT[2032*9 +: 8], 
          INIT[2031*9 +: 8], INIT[2030*9 +: 8], INIT[2029*9 +: 8], INIT[2028*9 +: 8], 
          INIT[2027*9 +: 8], INIT[2026*9 +: 8], INIT[2025*9 +: 8], INIT[2024*9 +: 8], 
          INIT[2023*9 +: 8], INIT[2022*9 +: 8], INIT[2021*9 +: 8], INIT[2020*9 +: 8], 
          INIT[2019*9 +: 8], INIT[2018*9 +: 8], INIT[2017*9 +: 8], INIT[2016*9 +: 8]}),
.INIT_40({INIT[2079*9 +: 8], INIT[2078*9 +: 8], INIT[2077*9 +: 8], INIT[2076*9 +: 8], 
          INIT[2075*9 +: 8], INIT[2074*9 +: 8], INIT[2073*9 +: 8], INIT[2072*9 +: 8], 
          INIT[2071*9 +: 8], INIT[2070*9 +: 8], INIT[2069*9 +: 8], INIT[2068*9 +: 8], 
          INIT[2067*9 +: 8], INIT[2066*9 +: 8], INIT[2065*9 +: 8], INIT[2064*9 +: 8], 
          INIT[2063*9 +: 8], INIT[2062*9 +: 8], INIT[2061*9 +: 8], INIT[2060*9 +: 8], 
          INIT[2059*9 +: 8], INIT[2058*9 +: 8], INIT[2057*9 +: 8], INIT[2056*9 +: 8], 
          INIT[2055*9 +: 8], INIT[2054*9 +: 8], INIT[2053*9 +: 8], INIT[2052*9 +: 8], 
          INIT[2051*9 +: 8], INIT[2050*9 +: 8], INIT[2049*9 +: 8], INIT[2048*9 +: 8]}),
.INIT_41({INIT[2111*9 +: 8], INIT[2110*9 +: 8], INIT[2109*9 +: 8], INIT[2108*9 +: 8], 
          INIT[2107*9 +: 8], INIT[2106*9 +: 8], INIT[2105*9 +: 8], INIT[2104*9 +: 8], 
          INIT[2103*9 +: 8], INIT[2102*9 +: 8], INIT[2101*9 +: 8], INIT[2100*9 +: 8], 
          INIT[2099*9 +: 8], INIT[2098*9 +: 8], INIT[2097*9 +: 8], INIT[2096*9 +: 8], 
          INIT[2095*9 +: 8], INIT[2094*9 +: 8], INIT[2093*9 +: 8], INIT[2092*9 +: 8], 
          INIT[2091*9 +: 8], INIT[2090*9 +: 8], INIT[2089*9 +: 8], INIT[2088*9 +: 8], 
          INIT[2087*9 +: 8], INIT[2086*9 +: 8], INIT[2085*9 +: 8], INIT[2084*9 +: 8], 
          INIT[2083*9 +: 8], INIT[2082*9 +: 8], INIT[2081*9 +: 8], INIT[2080*9 +: 8]}),
.INIT_42({INIT[2143*9 +: 8], INIT[2142*9 +: 8], INIT[2141*9 +: 8], INIT[2140*9 +: 8], 
          INIT[2139*9 +: 8], INIT[2138*9 +: 8], INIT[2137*9 +: 8], INIT[2136*9 +: 8], 
          INIT[2135*9 +: 8], INIT[2134*9 +: 8], INIT[2133*9 +: 8], INIT[2132*9 +: 8], 
          INIT[2131*9 +: 8], INIT[2130*9 +: 8], INIT[2129*9 +: 8], INIT[2128*9 +: 8], 
          INIT[2127*9 +: 8], INIT[2126*9 +: 8], INIT[2125*9 +: 8], INIT[2124*9 +: 8], 
          INIT[2123*9 +: 8], INIT[2122*9 +: 8], INIT[2121*9 +: 8], INIT[2120*9 +: 8], 
          INIT[2119*9 +: 8], INIT[2118*9 +: 8], INIT[2117*9 +: 8], INIT[2116*9 +: 8], 
          INIT[2115*9 +: 8], INIT[2114*9 +: 8], INIT[2113*9 +: 8], INIT[2112*9 +: 8]}),
.INIT_43({INIT[2175*9 +: 8], INIT[2174*9 +: 8], INIT[2173*9 +: 8], INIT[2172*9 +: 8], 
          INIT[2171*9 +: 8], INIT[2170*9 +: 8], INIT[2169*9 +: 8], INIT[2168*9 +: 8], 
          INIT[2167*9 +: 8], INIT[2166*9 +: 8], INIT[2165*9 +: 8], INIT[2164*9 +: 8], 
          INIT[2163*9 +: 8], INIT[2162*9 +: 8], INIT[2161*9 +: 8], INIT[2160*9 +: 8], 
          INIT[2159*9 +: 8], INIT[2158*9 +: 8], INIT[2157*9 +: 8], INIT[2156*9 +: 8], 
          INIT[2155*9 +: 8], INIT[2154*9 +: 8], INIT[2153*9 +: 8], INIT[2152*9 +: 8], 
          INIT[2151*9 +: 8], INIT[2150*9 +: 8], INIT[2149*9 +: 8], INIT[2148*9 +: 8], 
          INIT[2147*9 +: 8], INIT[2146*9 +: 8], INIT[2145*9 +: 8], INIT[2144*9 +: 8]}),
.INIT_44({INIT[2207*9 +: 8], INIT[2206*9 +: 8], INIT[2205*9 +: 8], INIT[2204*9 +: 8], 
          INIT[2203*9 +: 8], INIT[2202*9 +: 8], INIT[2201*9 +: 8], INIT[2200*9 +: 8], 
          INIT[2199*9 +: 8], INIT[2198*9 +: 8], INIT[2197*9 +: 8], INIT[2196*9 +: 8], 
          INIT[2195*9 +: 8], INIT[2194*9 +: 8], INIT[2193*9 +: 8], INIT[2192*9 +: 8], 
          INIT[2191*9 +: 8], INIT[2190*9 +: 8], INIT[2189*9 +: 8], INIT[2188*9 +: 8], 
          INIT[2187*9 +: 8], INIT[2186*9 +: 8], INIT[2185*9 +: 8], INIT[2184*9 +: 8], 
          INIT[2183*9 +: 8], INIT[2182*9 +: 8], INIT[2181*9 +: 8], INIT[2180*9 +: 8], 
          INIT[2179*9 +: 8], INIT[2178*9 +: 8], INIT[2177*9 +: 8], INIT[2176*9 +: 8]}),
.INIT_45({INIT[2239*9 +: 8], INIT[2238*9 +: 8], INIT[2237*9 +: 8], INIT[2236*9 +: 8], 
          INIT[2235*9 +: 8], INIT[2234*9 +: 8], INIT[2233*9 +: 8], INIT[2232*9 +: 8], 
          INIT[2231*9 +: 8], INIT[2230*9 +: 8], INIT[2229*9 +: 8], INIT[2228*9 +: 8], 
          INIT[2227*9 +: 8], INIT[2226*9 +: 8], INIT[2225*9 +: 8], INIT[2224*9 +: 8], 
          INIT[2223*9 +: 8], INIT[2222*9 +: 8], INIT[2221*9 +: 8], INIT[2220*9 +: 8], 
          INIT[2219*9 +: 8], INIT[2218*9 +: 8], INIT[2217*9 +: 8], INIT[2216*9 +: 8], 
          INIT[2215*9 +: 8], INIT[2214*9 +: 8], INIT[2213*9 +: 8], INIT[2212*9 +: 8], 
          INIT[2211*9 +: 8], INIT[2210*9 +: 8], INIT[2209*9 +: 8], INIT[2208*9 +: 8]}),
.INIT_46({INIT[2271*9 +: 8], INIT[2270*9 +: 8], INIT[2269*9 +: 8], INIT[2268*9 +: 8], 
          INIT[2267*9 +: 8], INIT[2266*9 +: 8], INIT[2265*9 +: 8], INIT[2264*9 +: 8], 
          INIT[2263*9 +: 8], INIT[2262*9 +: 8], INIT[2261*9 +: 8], INIT[2260*9 +: 8], 
          INIT[2259*9 +: 8], INIT[2258*9 +: 8], INIT[2257*9 +: 8], INIT[2256*9 +: 8], 
          INIT[2255*9 +: 8], INIT[2254*9 +: 8], INIT[2253*9 +: 8], INIT[2252*9 +: 8], 
          INIT[2251*9 +: 8], INIT[2250*9 +: 8], INIT[2249*9 +: 8], INIT[2248*9 +: 8], 
          INIT[2247*9 +: 8], INIT[2246*9 +: 8], INIT[2245*9 +: 8], INIT[2244*9 +: 8], 
          INIT[2243*9 +: 8], INIT[2242*9 +: 8], INIT[2241*9 +: 8], INIT[2240*9 +: 8]}),
.INIT_47({INIT[2303*9 +: 8], INIT[2302*9 +: 8], INIT[2301*9 +: 8], INIT[2300*9 +: 8], 
          INIT[2299*9 +: 8], INIT[2298*9 +: 8], INIT[2297*9 +: 8], INIT[2296*9 +: 8], 
          INIT[2295*9 +: 8], INIT[2294*9 +: 8], INIT[2293*9 +: 8], INIT[2292*9 +: 8], 
          INIT[2291*9 +: 8], INIT[2290*9 +: 8], INIT[2289*9 +: 8], INIT[2288*9 +: 8], 
          INIT[2287*9 +: 8], INIT[2286*9 +: 8], INIT[2285*9 +: 8], INIT[2284*9 +: 8], 
          INIT[2283*9 +: 8], INIT[2282*9 +: 8], INIT[2281*9 +: 8], INIT[2280*9 +: 8], 
          INIT[2279*9 +: 8], INIT[2278*9 +: 8], INIT[2277*9 +: 8], INIT[2276*9 +: 8], 
          INIT[2275*9 +: 8], INIT[2274*9 +: 8], INIT[2273*9 +: 8], INIT[2272*9 +: 8]}),
.INIT_48({INIT[2335*9 +: 8], INIT[2334*9 +: 8], INIT[2333*9 +: 8], INIT[2332*9 +: 8], 
          INIT[2331*9 +: 8], INIT[2330*9 +: 8], INIT[2329*9 +: 8], INIT[2328*9 +: 8], 
          INIT[2327*9 +: 8], INIT[2326*9 +: 8], INIT[2325*9 +: 8], INIT[2324*9 +: 8], 
          INIT[2323*9 +: 8], INIT[2322*9 +: 8], INIT[2321*9 +: 8], INIT[2320*9 +: 8], 
          INIT[2319*9 +: 8], INIT[2318*9 +: 8], INIT[2317*9 +: 8], INIT[2316*9 +: 8], 
          INIT[2315*9 +: 8], INIT[2314*9 +: 8], INIT[2313*9 +: 8], INIT[2312*9 +: 8], 
          INIT[2311*9 +: 8], INIT[2310*9 +: 8], INIT[2309*9 +: 8], INIT[2308*9 +: 8], 
          INIT[2307*9 +: 8], INIT[2306*9 +: 8], INIT[2305*9 +: 8], INIT[2304*9 +: 8]}),
.INIT_49({INIT[2367*9 +: 8], INIT[2366*9 +: 8], INIT[2365*9 +: 8], INIT[2364*9 +: 8], 
          INIT[2363*9 +: 8], INIT[2362*9 +: 8], INIT[2361*9 +: 8], INIT[2360*9 +: 8], 
          INIT[2359*9 +: 8], INIT[2358*9 +: 8], INIT[2357*9 +: 8], INIT[2356*9 +: 8], 
          INIT[2355*9 +: 8], INIT[2354*9 +: 8], INIT[2353*9 +: 8], INIT[2352*9 +: 8], 
          INIT[2351*9 +: 8], INIT[2350*9 +: 8], INIT[2349*9 +: 8], INIT[2348*9 +: 8], 
          INIT[2347*9 +: 8], INIT[2346*9 +: 8], INIT[2345*9 +: 8], INIT[2344*9 +: 8], 
          INIT[2343*9 +: 8], INIT[2342*9 +: 8], INIT[2341*9 +: 8], INIT[2340*9 +: 8], 
          INIT[2339*9 +: 8], INIT[2338*9 +: 8], INIT[2337*9 +: 8], INIT[2336*9 +: 8]}),
.INIT_4A({INIT[2399*9 +: 8], INIT[2398*9 +: 8], INIT[2397*9 +: 8], INIT[2396*9 +: 8], 
          INIT[2395*9 +: 8], INIT[2394*9 +: 8], INIT[2393*9 +: 8], INIT[2392*9 +: 8], 
          INIT[2391*9 +: 8], INIT[2390*9 +: 8], INIT[2389*9 +: 8], INIT[2388*9 +: 8], 
          INIT[2387*9 +: 8], INIT[2386*9 +: 8], INIT[2385*9 +: 8], INIT[2384*9 +: 8], 
          INIT[2383*9 +: 8], INIT[2382*9 +: 8], INIT[2381*9 +: 8], INIT[2380*9 +: 8], 
          INIT[2379*9 +: 8], INIT[2378*9 +: 8], INIT[2377*9 +: 8], INIT[2376*9 +: 8], 
          INIT[2375*9 +: 8], INIT[2374*9 +: 8], INIT[2373*9 +: 8], INIT[2372*9 +: 8], 
          INIT[2371*9 +: 8], INIT[2370*9 +: 8], INIT[2369*9 +: 8], INIT[2368*9 +: 8]}),
.INIT_4B({INIT[2431*9 +: 8], INIT[2430*9 +: 8], INIT[2429*9 +: 8], INIT[2428*9 +: 8], 
          INIT[2427*9 +: 8], INIT[2426*9 +: 8], INIT[2425*9 +: 8], INIT[2424*9 +: 8], 
          INIT[2423*9 +: 8], INIT[2422*9 +: 8], INIT[2421*9 +: 8], INIT[2420*9 +: 8], 
          INIT[2419*9 +: 8], INIT[2418*9 +: 8], INIT[2417*9 +: 8], INIT[2416*9 +: 8], 
          INIT[2415*9 +: 8], INIT[2414*9 +: 8], INIT[2413*9 +: 8], INIT[2412*9 +: 8], 
          INIT[2411*9 +: 8], INIT[2410*9 +: 8], INIT[2409*9 +: 8], INIT[2408*9 +: 8], 
          INIT[2407*9 +: 8], INIT[2406*9 +: 8], INIT[2405*9 +: 8], INIT[2404*9 +: 8], 
          INIT[2403*9 +: 8], INIT[2402*9 +: 8], INIT[2401*9 +: 8], INIT[2400*9 +: 8]}),
.INIT_4C({INIT[2463*9 +: 8], INIT[2462*9 +: 8], INIT[2461*9 +: 8], INIT[2460*9 +: 8], 
          INIT[2459*9 +: 8], INIT[2458*9 +: 8], INIT[2457*9 +: 8], INIT[2456*9 +: 8], 
          INIT[2455*9 +: 8], INIT[2454*9 +: 8], INIT[2453*9 +: 8], INIT[2452*9 +: 8], 
          INIT[2451*9 +: 8], INIT[2450*9 +: 8], INIT[2449*9 +: 8], INIT[2448*9 +: 8], 
          INIT[2447*9 +: 8], INIT[2446*9 +: 8], INIT[2445*9 +: 8], INIT[2444*9 +: 8], 
          INIT[2443*9 +: 8], INIT[2442*9 +: 8], INIT[2441*9 +: 8], INIT[2440*9 +: 8], 
          INIT[2439*9 +: 8], INIT[2438*9 +: 8], INIT[2437*9 +: 8], INIT[2436*9 +: 8], 
          INIT[2435*9 +: 8], INIT[2434*9 +: 8], INIT[2433*9 +: 8], INIT[2432*9 +: 8]}),
.INIT_4D({INIT[2495*9 +: 8], INIT[2494*9 +: 8], INIT[2493*9 +: 8], INIT[2492*9 +: 8], 
          INIT[2491*9 +: 8], INIT[2490*9 +: 8], INIT[2489*9 +: 8], INIT[2488*9 +: 8], 
          INIT[2487*9 +: 8], INIT[2486*9 +: 8], INIT[2485*9 +: 8], INIT[2484*9 +: 8], 
          INIT[2483*9 +: 8], INIT[2482*9 +: 8], INIT[2481*9 +: 8], INIT[2480*9 +: 8], 
          INIT[2479*9 +: 8], INIT[2478*9 +: 8], INIT[2477*9 +: 8], INIT[2476*9 +: 8], 
          INIT[2475*9 +: 8], INIT[2474*9 +: 8], INIT[2473*9 +: 8], INIT[2472*9 +: 8], 
          INIT[2471*9 +: 8], INIT[2470*9 +: 8], INIT[2469*9 +: 8], INIT[2468*9 +: 8], 
          INIT[2467*9 +: 8], INIT[2466*9 +: 8], INIT[2465*9 +: 8], INIT[2464*9 +: 8]}),
.INIT_4E({INIT[2527*9 +: 8], INIT[2526*9 +: 8], INIT[2525*9 +: 8], INIT[2524*9 +: 8], 
          INIT[2523*9 +: 8], INIT[2522*9 +: 8], INIT[2521*9 +: 8], INIT[2520*9 +: 8], 
          INIT[2519*9 +: 8], INIT[2518*9 +: 8], INIT[2517*9 +: 8], INIT[2516*9 +: 8], 
          INIT[2515*9 +: 8], INIT[2514*9 +: 8], INIT[2513*9 +: 8], INIT[2512*9 +: 8], 
          INIT[2511*9 +: 8], INIT[2510*9 +: 8], INIT[2509*9 +: 8], INIT[2508*9 +: 8], 
          INIT[2507*9 +: 8], INIT[2506*9 +: 8], INIT[2505*9 +: 8], INIT[2504*9 +: 8], 
          INIT[2503*9 +: 8], INIT[2502*9 +: 8], INIT[2501*9 +: 8], INIT[2500*9 +: 8], 
          INIT[2499*9 +: 8], INIT[2498*9 +: 8], INIT[2497*9 +: 8], INIT[2496*9 +: 8]}),
.INIT_4F({INIT[2559*9 +: 8], INIT[2558*9 +: 8], INIT[2557*9 +: 8], INIT[2556*9 +: 8], 
          INIT[2555*9 +: 8], INIT[2554*9 +: 8], INIT[2553*9 +: 8], INIT[2552*9 +: 8], 
          INIT[2551*9 +: 8], INIT[2550*9 +: 8], INIT[2549*9 +: 8], INIT[2548*9 +: 8], 
          INIT[2547*9 +: 8], INIT[2546*9 +: 8], INIT[2545*9 +: 8], INIT[2544*9 +: 8], 
          INIT[2543*9 +: 8], INIT[2542*9 +: 8], INIT[2541*9 +: 8], INIT[2540*9 +: 8], 
          INIT[2539*9 +: 8], INIT[2538*9 +: 8], INIT[2537*9 +: 8], INIT[2536*9 +: 8], 
          INIT[2535*9 +: 8], INIT[2534*9 +: 8], INIT[2533*9 +: 8], INIT[2532*9 +: 8], 
          INIT[2531*9 +: 8], INIT[2530*9 +: 8], INIT[2529*9 +: 8], INIT[2528*9 +: 8]}),
.INIT_50({INIT[2591*9 +: 8], INIT[2590*9 +: 8], INIT[2589*9 +: 8], INIT[2588*9 +: 8], 
          INIT[2587*9 +: 8], INIT[2586*9 +: 8], INIT[2585*9 +: 8], INIT[2584*9 +: 8], 
          INIT[2583*9 +: 8], INIT[2582*9 +: 8], INIT[2581*9 +: 8], INIT[2580*9 +: 8], 
          INIT[2579*9 +: 8], INIT[2578*9 +: 8], INIT[2577*9 +: 8], INIT[2576*9 +: 8], 
          INIT[2575*9 +: 8], INIT[2574*9 +: 8], INIT[2573*9 +: 8], INIT[2572*9 +: 8], 
          INIT[2571*9 +: 8], INIT[2570*9 +: 8], INIT[2569*9 +: 8], INIT[2568*9 +: 8], 
          INIT[2567*9 +: 8], INIT[2566*9 +: 8], INIT[2565*9 +: 8], INIT[2564*9 +: 8], 
          INIT[2563*9 +: 8], INIT[2562*9 +: 8], INIT[2561*9 +: 8], INIT[2560*9 +: 8]}),
.INIT_51({INIT[2623*9 +: 8], INIT[2622*9 +: 8], INIT[2621*9 +: 8], INIT[2620*9 +: 8], 
          INIT[2619*9 +: 8], INIT[2618*9 +: 8], INIT[2617*9 +: 8], INIT[2616*9 +: 8], 
          INIT[2615*9 +: 8], INIT[2614*9 +: 8], INIT[2613*9 +: 8], INIT[2612*9 +: 8], 
          INIT[2611*9 +: 8], INIT[2610*9 +: 8], INIT[2609*9 +: 8], INIT[2608*9 +: 8], 
          INIT[2607*9 +: 8], INIT[2606*9 +: 8], INIT[2605*9 +: 8], INIT[2604*9 +: 8], 
          INIT[2603*9 +: 8], INIT[2602*9 +: 8], INIT[2601*9 +: 8], INIT[2600*9 +: 8], 
          INIT[2599*9 +: 8], INIT[2598*9 +: 8], INIT[2597*9 +: 8], INIT[2596*9 +: 8], 
          INIT[2595*9 +: 8], INIT[2594*9 +: 8], INIT[2593*9 +: 8], INIT[2592*9 +: 8]}),
.INIT_52({INIT[2655*9 +: 8], INIT[2654*9 +: 8], INIT[2653*9 +: 8], INIT[2652*9 +: 8], 
          INIT[2651*9 +: 8], INIT[2650*9 +: 8], INIT[2649*9 +: 8], INIT[2648*9 +: 8], 
          INIT[2647*9 +: 8], INIT[2646*9 +: 8], INIT[2645*9 +: 8], INIT[2644*9 +: 8], 
          INIT[2643*9 +: 8], INIT[2642*9 +: 8], INIT[2641*9 +: 8], INIT[2640*9 +: 8], 
          INIT[2639*9 +: 8], INIT[2638*9 +: 8], INIT[2637*9 +: 8], INIT[2636*9 +: 8], 
          INIT[2635*9 +: 8], INIT[2634*9 +: 8], INIT[2633*9 +: 8], INIT[2632*9 +: 8], 
          INIT[2631*9 +: 8], INIT[2630*9 +: 8], INIT[2629*9 +: 8], INIT[2628*9 +: 8], 
          INIT[2627*9 +: 8], INIT[2626*9 +: 8], INIT[2625*9 +: 8], INIT[2624*9 +: 8]}),
.INIT_53({INIT[2687*9 +: 8], INIT[2686*9 +: 8], INIT[2685*9 +: 8], INIT[2684*9 +: 8], 
          INIT[2683*9 +: 8], INIT[2682*9 +: 8], INIT[2681*9 +: 8], INIT[2680*9 +: 8], 
          INIT[2679*9 +: 8], INIT[2678*9 +: 8], INIT[2677*9 +: 8], INIT[2676*9 +: 8], 
          INIT[2675*9 +: 8], INIT[2674*9 +: 8], INIT[2673*9 +: 8], INIT[2672*9 +: 8], 
          INIT[2671*9 +: 8], INIT[2670*9 +: 8], INIT[2669*9 +: 8], INIT[2668*9 +: 8], 
          INIT[2667*9 +: 8], INIT[2666*9 +: 8], INIT[2665*9 +: 8], INIT[2664*9 +: 8], 
          INIT[2663*9 +: 8], INIT[2662*9 +: 8], INIT[2661*9 +: 8], INIT[2660*9 +: 8], 
          INIT[2659*9 +: 8], INIT[2658*9 +: 8], INIT[2657*9 +: 8], INIT[2656*9 +: 8]}),
.INIT_54({INIT[2719*9 +: 8], INIT[2718*9 +: 8], INIT[2717*9 +: 8], INIT[2716*9 +: 8], 
          INIT[2715*9 +: 8], INIT[2714*9 +: 8], INIT[2713*9 +: 8], INIT[2712*9 +: 8], 
          INIT[2711*9 +: 8], INIT[2710*9 +: 8], INIT[2709*9 +: 8], INIT[2708*9 +: 8], 
          INIT[2707*9 +: 8], INIT[2706*9 +: 8], INIT[2705*9 +: 8], INIT[2704*9 +: 8], 
          INIT[2703*9 +: 8], INIT[2702*9 +: 8], INIT[2701*9 +: 8], INIT[2700*9 +: 8], 
          INIT[2699*9 +: 8], INIT[2698*9 +: 8], INIT[2697*9 +: 8], INIT[2696*9 +: 8], 
          INIT[2695*9 +: 8], INIT[2694*9 +: 8], INIT[2693*9 +: 8], INIT[2692*9 +: 8], 
          INIT[2691*9 +: 8], INIT[2690*9 +: 8], INIT[2689*9 +: 8], INIT[2688*9 +: 8]}),
.INIT_55({INIT[2751*9 +: 8], INIT[2750*9 +: 8], INIT[2749*9 +: 8], INIT[2748*9 +: 8], 
          INIT[2747*9 +: 8], INIT[2746*9 +: 8], INIT[2745*9 +: 8], INIT[2744*9 +: 8], 
          INIT[2743*9 +: 8], INIT[2742*9 +: 8], INIT[2741*9 +: 8], INIT[2740*9 +: 8], 
          INIT[2739*9 +: 8], INIT[2738*9 +: 8], INIT[2737*9 +: 8], INIT[2736*9 +: 8], 
          INIT[2735*9 +: 8], INIT[2734*9 +: 8], INIT[2733*9 +: 8], INIT[2732*9 +: 8], 
          INIT[2731*9 +: 8], INIT[2730*9 +: 8], INIT[2729*9 +: 8], INIT[2728*9 +: 8], 
          INIT[2727*9 +: 8], INIT[2726*9 +: 8], INIT[2725*9 +: 8], INIT[2724*9 +: 8], 
          INIT[2723*9 +: 8], INIT[2722*9 +: 8], INIT[2721*9 +: 8], INIT[2720*9 +: 8]}),
.INIT_56({INIT[2783*9 +: 8], INIT[2782*9 +: 8], INIT[2781*9 +: 8], INIT[2780*9 +: 8], 
          INIT[2779*9 +: 8], INIT[2778*9 +: 8], INIT[2777*9 +: 8], INIT[2776*9 +: 8], 
          INIT[2775*9 +: 8], INIT[2774*9 +: 8], INIT[2773*9 +: 8], INIT[2772*9 +: 8], 
          INIT[2771*9 +: 8], INIT[2770*9 +: 8], INIT[2769*9 +: 8], INIT[2768*9 +: 8], 
          INIT[2767*9 +: 8], INIT[2766*9 +: 8], INIT[2765*9 +: 8], INIT[2764*9 +: 8], 
          INIT[2763*9 +: 8], INIT[2762*9 +: 8], INIT[2761*9 +: 8], INIT[2760*9 +: 8], 
          INIT[2759*9 +: 8], INIT[2758*9 +: 8], INIT[2757*9 +: 8], INIT[2756*9 +: 8], 
          INIT[2755*9 +: 8], INIT[2754*9 +: 8], INIT[2753*9 +: 8], INIT[2752*9 +: 8]}),
.INIT_57({INIT[2815*9 +: 8], INIT[2814*9 +: 8], INIT[2813*9 +: 8], INIT[2812*9 +: 8], 
          INIT[2811*9 +: 8], INIT[2810*9 +: 8], INIT[2809*9 +: 8], INIT[2808*9 +: 8], 
          INIT[2807*9 +: 8], INIT[2806*9 +: 8], INIT[2805*9 +: 8], INIT[2804*9 +: 8], 
          INIT[2803*9 +: 8], INIT[2802*9 +: 8], INIT[2801*9 +: 8], INIT[2800*9 +: 8], 
          INIT[2799*9 +: 8], INIT[2798*9 +: 8], INIT[2797*9 +: 8], INIT[2796*9 +: 8], 
          INIT[2795*9 +: 8], INIT[2794*9 +: 8], INIT[2793*9 +: 8], INIT[2792*9 +: 8], 
          INIT[2791*9 +: 8], INIT[2790*9 +: 8], INIT[2789*9 +: 8], INIT[2788*9 +: 8], 
          INIT[2787*9 +: 8], INIT[2786*9 +: 8], INIT[2785*9 +: 8], INIT[2784*9 +: 8]}),
.INIT_58({INIT[2847*9 +: 8], INIT[2846*9 +: 8], INIT[2845*9 +: 8], INIT[2844*9 +: 8], 
          INIT[2843*9 +: 8], INIT[2842*9 +: 8], INIT[2841*9 +: 8], INIT[2840*9 +: 8], 
          INIT[2839*9 +: 8], INIT[2838*9 +: 8], INIT[2837*9 +: 8], INIT[2836*9 +: 8], 
          INIT[2835*9 +: 8], INIT[2834*9 +: 8], INIT[2833*9 +: 8], INIT[2832*9 +: 8], 
          INIT[2831*9 +: 8], INIT[2830*9 +: 8], INIT[2829*9 +: 8], INIT[2828*9 +: 8], 
          INIT[2827*9 +: 8], INIT[2826*9 +: 8], INIT[2825*9 +: 8], INIT[2824*9 +: 8], 
          INIT[2823*9 +: 8], INIT[2822*9 +: 8], INIT[2821*9 +: 8], INIT[2820*9 +: 8], 
          INIT[2819*9 +: 8], INIT[2818*9 +: 8], INIT[2817*9 +: 8], INIT[2816*9 +: 8]}),
.INIT_59({INIT[2879*9 +: 8], INIT[2878*9 +: 8], INIT[2877*9 +: 8], INIT[2876*9 +: 8], 
          INIT[2875*9 +: 8], INIT[2874*9 +: 8], INIT[2873*9 +: 8], INIT[2872*9 +: 8], 
          INIT[2871*9 +: 8], INIT[2870*9 +: 8], INIT[2869*9 +: 8], INIT[2868*9 +: 8], 
          INIT[2867*9 +: 8], INIT[2866*9 +: 8], INIT[2865*9 +: 8], INIT[2864*9 +: 8], 
          INIT[2863*9 +: 8], INIT[2862*9 +: 8], INIT[2861*9 +: 8], INIT[2860*9 +: 8], 
          INIT[2859*9 +: 8], INIT[2858*9 +: 8], INIT[2857*9 +: 8], INIT[2856*9 +: 8], 
          INIT[2855*9 +: 8], INIT[2854*9 +: 8], INIT[2853*9 +: 8], INIT[2852*9 +: 8], 
          INIT[2851*9 +: 8], INIT[2850*9 +: 8], INIT[2849*9 +: 8], INIT[2848*9 +: 8]}),
.INIT_5A({INIT[2911*9 +: 8], INIT[2910*9 +: 8], INIT[2909*9 +: 8], INIT[2908*9 +: 8], 
          INIT[2907*9 +: 8], INIT[2906*9 +: 8], INIT[2905*9 +: 8], INIT[2904*9 +: 8], 
          INIT[2903*9 +: 8], INIT[2902*9 +: 8], INIT[2901*9 +: 8], INIT[2900*9 +: 8], 
          INIT[2899*9 +: 8], INIT[2898*9 +: 8], INIT[2897*9 +: 8], INIT[2896*9 +: 8], 
          INIT[2895*9 +: 8], INIT[2894*9 +: 8], INIT[2893*9 +: 8], INIT[2892*9 +: 8], 
          INIT[2891*9 +: 8], INIT[2890*9 +: 8], INIT[2889*9 +: 8], INIT[2888*9 +: 8], 
          INIT[2887*9 +: 8], INIT[2886*9 +: 8], INIT[2885*9 +: 8], INIT[2884*9 +: 8], 
          INIT[2883*9 +: 8], INIT[2882*9 +: 8], INIT[2881*9 +: 8], INIT[2880*9 +: 8]}),
.INIT_5B({INIT[2943*9 +: 8], INIT[2942*9 +: 8], INIT[2941*9 +: 8], INIT[2940*9 +: 8], 
          INIT[2939*9 +: 8], INIT[2938*9 +: 8], INIT[2937*9 +: 8], INIT[2936*9 +: 8], 
          INIT[2935*9 +: 8], INIT[2934*9 +: 8], INIT[2933*9 +: 8], INIT[2932*9 +: 8], 
          INIT[2931*9 +: 8], INIT[2930*9 +: 8], INIT[2929*9 +: 8], INIT[2928*9 +: 8], 
          INIT[2927*9 +: 8], INIT[2926*9 +: 8], INIT[2925*9 +: 8], INIT[2924*9 +: 8], 
          INIT[2923*9 +: 8], INIT[2922*9 +: 8], INIT[2921*9 +: 8], INIT[2920*9 +: 8], 
          INIT[2919*9 +: 8], INIT[2918*9 +: 8], INIT[2917*9 +: 8], INIT[2916*9 +: 8], 
          INIT[2915*9 +: 8], INIT[2914*9 +: 8], INIT[2913*9 +: 8], INIT[2912*9 +: 8]}),
.INIT_5C({INIT[2975*9 +: 8], INIT[2974*9 +: 8], INIT[2973*9 +: 8], INIT[2972*9 +: 8], 
          INIT[2971*9 +: 8], INIT[2970*9 +: 8], INIT[2969*9 +: 8], INIT[2968*9 +: 8], 
          INIT[2967*9 +: 8], INIT[2966*9 +: 8], INIT[2965*9 +: 8], INIT[2964*9 +: 8], 
          INIT[2963*9 +: 8], INIT[2962*9 +: 8], INIT[2961*9 +: 8], INIT[2960*9 +: 8], 
          INIT[2959*9 +: 8], INIT[2958*9 +: 8], INIT[2957*9 +: 8], INIT[2956*9 +: 8], 
          INIT[2955*9 +: 8], INIT[2954*9 +: 8], INIT[2953*9 +: 8], INIT[2952*9 +: 8], 
          INIT[2951*9 +: 8], INIT[2950*9 +: 8], INIT[2949*9 +: 8], INIT[2948*9 +: 8], 
          INIT[2947*9 +: 8], INIT[2946*9 +: 8], INIT[2945*9 +: 8], INIT[2944*9 +: 8]}),
.INIT_5D({INIT[3007*9 +: 8], INIT[3006*9 +: 8], INIT[3005*9 +: 8], INIT[3004*9 +: 8], 
          INIT[3003*9 +: 8], INIT[3002*9 +: 8], INIT[3001*9 +: 8], INIT[3000*9 +: 8], 
          INIT[2999*9 +: 8], INIT[2998*9 +: 8], INIT[2997*9 +: 8], INIT[2996*9 +: 8], 
          INIT[2995*9 +: 8], INIT[2994*9 +: 8], INIT[2993*9 +: 8], INIT[2992*9 +: 8], 
          INIT[2991*9 +: 8], INIT[2990*9 +: 8], INIT[2989*9 +: 8], INIT[2988*9 +: 8], 
          INIT[2987*9 +: 8], INIT[2986*9 +: 8], INIT[2985*9 +: 8], INIT[2984*9 +: 8], 
          INIT[2983*9 +: 8], INIT[2982*9 +: 8], INIT[2981*9 +: 8], INIT[2980*9 +: 8], 
          INIT[2979*9 +: 8], INIT[2978*9 +: 8], INIT[2977*9 +: 8], INIT[2976*9 +: 8]}),
.INIT_5E({INIT[3039*9 +: 8], INIT[3038*9 +: 8], INIT[3037*9 +: 8], INIT[3036*9 +: 8], 
          INIT[3035*9 +: 8], INIT[3034*9 +: 8], INIT[3033*9 +: 8], INIT[3032*9 +: 8], 
          INIT[3031*9 +: 8], INIT[3030*9 +: 8], INIT[3029*9 +: 8], INIT[3028*9 +: 8], 
          INIT[3027*9 +: 8], INIT[3026*9 +: 8], INIT[3025*9 +: 8], INIT[3024*9 +: 8], 
          INIT[3023*9 +: 8], INIT[3022*9 +: 8], INIT[3021*9 +: 8], INIT[3020*9 +: 8], 
          INIT[3019*9 +: 8], INIT[3018*9 +: 8], INIT[3017*9 +: 8], INIT[3016*9 +: 8], 
          INIT[3015*9 +: 8], INIT[3014*9 +: 8], INIT[3013*9 +: 8], INIT[3012*9 +: 8], 
          INIT[3011*9 +: 8], INIT[3010*9 +: 8], INIT[3009*9 +: 8], INIT[3008*9 +: 8]}),
.INIT_5F({INIT[3071*9 +: 8], INIT[3070*9 +: 8], INIT[3069*9 +: 8], INIT[3068*9 +: 8], 
          INIT[3067*9 +: 8], INIT[3066*9 +: 8], INIT[3065*9 +: 8], INIT[3064*9 +: 8], 
          INIT[3063*9 +: 8], INIT[3062*9 +: 8], INIT[3061*9 +: 8], INIT[3060*9 +: 8], 
          INIT[3059*9 +: 8], INIT[3058*9 +: 8], INIT[3057*9 +: 8], INIT[3056*9 +: 8], 
          INIT[3055*9 +: 8], INIT[3054*9 +: 8], INIT[3053*9 +: 8], INIT[3052*9 +: 8], 
          INIT[3051*9 +: 8], INIT[3050*9 +: 8], INIT[3049*9 +: 8], INIT[3048*9 +: 8], 
          INIT[3047*9 +: 8], INIT[3046*9 +: 8], INIT[3045*9 +: 8], INIT[3044*9 +: 8], 
          INIT[3043*9 +: 8], INIT[3042*9 +: 8], INIT[3041*9 +: 8], INIT[3040*9 +: 8]}),
.INIT_60({INIT[3103*9 +: 8], INIT[3102*9 +: 8], INIT[3101*9 +: 8], INIT[3100*9 +: 8], 
          INIT[3099*9 +: 8], INIT[3098*9 +: 8], INIT[3097*9 +: 8], INIT[3096*9 +: 8], 
          INIT[3095*9 +: 8], INIT[3094*9 +: 8], INIT[3093*9 +: 8], INIT[3092*9 +: 8], 
          INIT[3091*9 +: 8], INIT[3090*9 +: 8], INIT[3089*9 +: 8], INIT[3088*9 +: 8], 
          INIT[3087*9 +: 8], INIT[3086*9 +: 8], INIT[3085*9 +: 8], INIT[3084*9 +: 8], 
          INIT[3083*9 +: 8], INIT[3082*9 +: 8], INIT[3081*9 +: 8], INIT[3080*9 +: 8], 
          INIT[3079*9 +: 8], INIT[3078*9 +: 8], INIT[3077*9 +: 8], INIT[3076*9 +: 8], 
          INIT[3075*9 +: 8], INIT[3074*9 +: 8], INIT[3073*9 +: 8], INIT[3072*9 +: 8]}),
.INIT_61({INIT[3135*9 +: 8], INIT[3134*9 +: 8], INIT[3133*9 +: 8], INIT[3132*9 +: 8], 
          INIT[3131*9 +: 8], INIT[3130*9 +: 8], INIT[3129*9 +: 8], INIT[3128*9 +: 8], 
          INIT[3127*9 +: 8], INIT[3126*9 +: 8], INIT[3125*9 +: 8], INIT[3124*9 +: 8], 
          INIT[3123*9 +: 8], INIT[3122*9 +: 8], INIT[3121*9 +: 8], INIT[3120*9 +: 8], 
          INIT[3119*9 +: 8], INIT[3118*9 +: 8], INIT[3117*9 +: 8], INIT[3116*9 +: 8], 
          INIT[3115*9 +: 8], INIT[3114*9 +: 8], INIT[3113*9 +: 8], INIT[3112*9 +: 8], 
          INIT[3111*9 +: 8], INIT[3110*9 +: 8], INIT[3109*9 +: 8], INIT[3108*9 +: 8], 
          INIT[3107*9 +: 8], INIT[3106*9 +: 8], INIT[3105*9 +: 8], INIT[3104*9 +: 8]}),
.INIT_62({INIT[3167*9 +: 8], INIT[3166*9 +: 8], INIT[3165*9 +: 8], INIT[3164*9 +: 8], 
          INIT[3163*9 +: 8], INIT[3162*9 +: 8], INIT[3161*9 +: 8], INIT[3160*9 +: 8], 
          INIT[3159*9 +: 8], INIT[3158*9 +: 8], INIT[3157*9 +: 8], INIT[3156*9 +: 8], 
          INIT[3155*9 +: 8], INIT[3154*9 +: 8], INIT[3153*9 +: 8], INIT[3152*9 +: 8], 
          INIT[3151*9 +: 8], INIT[3150*9 +: 8], INIT[3149*9 +: 8], INIT[3148*9 +: 8], 
          INIT[3147*9 +: 8], INIT[3146*9 +: 8], INIT[3145*9 +: 8], INIT[3144*9 +: 8], 
          INIT[3143*9 +: 8], INIT[3142*9 +: 8], INIT[3141*9 +: 8], INIT[3140*9 +: 8], 
          INIT[3139*9 +: 8], INIT[3138*9 +: 8], INIT[3137*9 +: 8], INIT[3136*9 +: 8]}),
.INIT_63({INIT[3199*9 +: 8], INIT[3198*9 +: 8], INIT[3197*9 +: 8], INIT[3196*9 +: 8], 
          INIT[3195*9 +: 8], INIT[3194*9 +: 8], INIT[3193*9 +: 8], INIT[3192*9 +: 8], 
          INIT[3191*9 +: 8], INIT[3190*9 +: 8], INIT[3189*9 +: 8], INIT[3188*9 +: 8], 
          INIT[3187*9 +: 8], INIT[3186*9 +: 8], INIT[3185*9 +: 8], INIT[3184*9 +: 8], 
          INIT[3183*9 +: 8], INIT[3182*9 +: 8], INIT[3181*9 +: 8], INIT[3180*9 +: 8], 
          INIT[3179*9 +: 8], INIT[3178*9 +: 8], INIT[3177*9 +: 8], INIT[3176*9 +: 8], 
          INIT[3175*9 +: 8], INIT[3174*9 +: 8], INIT[3173*9 +: 8], INIT[3172*9 +: 8], 
          INIT[3171*9 +: 8], INIT[3170*9 +: 8], INIT[3169*9 +: 8], INIT[3168*9 +: 8]}),
.INIT_64({INIT[3231*9 +: 8], INIT[3230*9 +: 8], INIT[3229*9 +: 8], INIT[3228*9 +: 8], 
          INIT[3227*9 +: 8], INIT[3226*9 +: 8], INIT[3225*9 +: 8], INIT[3224*9 +: 8], 
          INIT[3223*9 +: 8], INIT[3222*9 +: 8], INIT[3221*9 +: 8], INIT[3220*9 +: 8], 
          INIT[3219*9 +: 8], INIT[3218*9 +: 8], INIT[3217*9 +: 8], INIT[3216*9 +: 8], 
          INIT[3215*9 +: 8], INIT[3214*9 +: 8], INIT[3213*9 +: 8], INIT[3212*9 +: 8], 
          INIT[3211*9 +: 8], INIT[3210*9 +: 8], INIT[3209*9 +: 8], INIT[3208*9 +: 8], 
          INIT[3207*9 +: 8], INIT[3206*9 +: 8], INIT[3205*9 +: 8], INIT[3204*9 +: 8], 
          INIT[3203*9 +: 8], INIT[3202*9 +: 8], INIT[3201*9 +: 8], INIT[3200*9 +: 8]}),
.INIT_65({INIT[3263*9 +: 8], INIT[3262*9 +: 8], INIT[3261*9 +: 8], INIT[3260*9 +: 8], 
          INIT[3259*9 +: 8], INIT[3258*9 +: 8], INIT[3257*9 +: 8], INIT[3256*9 +: 8], 
          INIT[3255*9 +: 8], INIT[3254*9 +: 8], INIT[3253*9 +: 8], INIT[3252*9 +: 8], 
          INIT[3251*9 +: 8], INIT[3250*9 +: 8], INIT[3249*9 +: 8], INIT[3248*9 +: 8], 
          INIT[3247*9 +: 8], INIT[3246*9 +: 8], INIT[3245*9 +: 8], INIT[3244*9 +: 8], 
          INIT[3243*9 +: 8], INIT[3242*9 +: 8], INIT[3241*9 +: 8], INIT[3240*9 +: 8], 
          INIT[3239*9 +: 8], INIT[3238*9 +: 8], INIT[3237*9 +: 8], INIT[3236*9 +: 8], 
          INIT[3235*9 +: 8], INIT[3234*9 +: 8], INIT[3233*9 +: 8], INIT[3232*9 +: 8]}),
.INIT_66({INIT[3295*9 +: 8], INIT[3294*9 +: 8], INIT[3293*9 +: 8], INIT[3292*9 +: 8], 
          INIT[3291*9 +: 8], INIT[3290*9 +: 8], INIT[3289*9 +: 8], INIT[3288*9 +: 8], 
          INIT[3287*9 +: 8], INIT[3286*9 +: 8], INIT[3285*9 +: 8], INIT[3284*9 +: 8], 
          INIT[3283*9 +: 8], INIT[3282*9 +: 8], INIT[3281*9 +: 8], INIT[3280*9 +: 8], 
          INIT[3279*9 +: 8], INIT[3278*9 +: 8], INIT[3277*9 +: 8], INIT[3276*9 +: 8], 
          INIT[3275*9 +: 8], INIT[3274*9 +: 8], INIT[3273*9 +: 8], INIT[3272*9 +: 8], 
          INIT[3271*9 +: 8], INIT[3270*9 +: 8], INIT[3269*9 +: 8], INIT[3268*9 +: 8], 
          INIT[3267*9 +: 8], INIT[3266*9 +: 8], INIT[3265*9 +: 8], INIT[3264*9 +: 8]}),
.INIT_67({INIT[3327*9 +: 8], INIT[3326*9 +: 8], INIT[3325*9 +: 8], INIT[3324*9 +: 8], 
          INIT[3323*9 +: 8], INIT[3322*9 +: 8], INIT[3321*9 +: 8], INIT[3320*9 +: 8], 
          INIT[3319*9 +: 8], INIT[3318*9 +: 8], INIT[3317*9 +: 8], INIT[3316*9 +: 8], 
          INIT[3315*9 +: 8], INIT[3314*9 +: 8], INIT[3313*9 +: 8], INIT[3312*9 +: 8], 
          INIT[3311*9 +: 8], INIT[3310*9 +: 8], INIT[3309*9 +: 8], INIT[3308*9 +: 8], 
          INIT[3307*9 +: 8], INIT[3306*9 +: 8], INIT[3305*9 +: 8], INIT[3304*9 +: 8], 
          INIT[3303*9 +: 8], INIT[3302*9 +: 8], INIT[3301*9 +: 8], INIT[3300*9 +: 8], 
          INIT[3299*9 +: 8], INIT[3298*9 +: 8], INIT[3297*9 +: 8], INIT[3296*9 +: 8]}),
.INIT_68({INIT[3359*9 +: 8], INIT[3358*9 +: 8], INIT[3357*9 +: 8], INIT[3356*9 +: 8], 
          INIT[3355*9 +: 8], INIT[3354*9 +: 8], INIT[3353*9 +: 8], INIT[3352*9 +: 8], 
          INIT[3351*9 +: 8], INIT[3350*9 +: 8], INIT[3349*9 +: 8], INIT[3348*9 +: 8], 
          INIT[3347*9 +: 8], INIT[3346*9 +: 8], INIT[3345*9 +: 8], INIT[3344*9 +: 8], 
          INIT[3343*9 +: 8], INIT[3342*9 +: 8], INIT[3341*9 +: 8], INIT[3340*9 +: 8], 
          INIT[3339*9 +: 8], INIT[3338*9 +: 8], INIT[3337*9 +: 8], INIT[3336*9 +: 8], 
          INIT[3335*9 +: 8], INIT[3334*9 +: 8], INIT[3333*9 +: 8], INIT[3332*9 +: 8], 
          INIT[3331*9 +: 8], INIT[3330*9 +: 8], INIT[3329*9 +: 8], INIT[3328*9 +: 8]}),
.INIT_69({INIT[3391*9 +: 8], INIT[3390*9 +: 8], INIT[3389*9 +: 8], INIT[3388*9 +: 8], 
          INIT[3387*9 +: 8], INIT[3386*9 +: 8], INIT[3385*9 +: 8], INIT[3384*9 +: 8], 
          INIT[3383*9 +: 8], INIT[3382*9 +: 8], INIT[3381*9 +: 8], INIT[3380*9 +: 8], 
          INIT[3379*9 +: 8], INIT[3378*9 +: 8], INIT[3377*9 +: 8], INIT[3376*9 +: 8], 
          INIT[3375*9 +: 8], INIT[3374*9 +: 8], INIT[3373*9 +: 8], INIT[3372*9 +: 8], 
          INIT[3371*9 +: 8], INIT[3370*9 +: 8], INIT[3369*9 +: 8], INIT[3368*9 +: 8], 
          INIT[3367*9 +: 8], INIT[3366*9 +: 8], INIT[3365*9 +: 8], INIT[3364*9 +: 8], 
          INIT[3363*9 +: 8], INIT[3362*9 +: 8], INIT[3361*9 +: 8], INIT[3360*9 +: 8]}),
.INIT_6A({INIT[3423*9 +: 8], INIT[3422*9 +: 8], INIT[3421*9 +: 8], INIT[3420*9 +: 8], 
          INIT[3419*9 +: 8], INIT[3418*9 +: 8], INIT[3417*9 +: 8], INIT[3416*9 +: 8], 
          INIT[3415*9 +: 8], INIT[3414*9 +: 8], INIT[3413*9 +: 8], INIT[3412*9 +: 8], 
          INIT[3411*9 +: 8], INIT[3410*9 +: 8], INIT[3409*9 +: 8], INIT[3408*9 +: 8], 
          INIT[3407*9 +: 8], INIT[3406*9 +: 8], INIT[3405*9 +: 8], INIT[3404*9 +: 8], 
          INIT[3403*9 +: 8], INIT[3402*9 +: 8], INIT[3401*9 +: 8], INIT[3400*9 +: 8], 
          INIT[3399*9 +: 8], INIT[3398*9 +: 8], INIT[3397*9 +: 8], INIT[3396*9 +: 8], 
          INIT[3395*9 +: 8], INIT[3394*9 +: 8], INIT[3393*9 +: 8], INIT[3392*9 +: 8]}),
.INIT_6B({INIT[3455*9 +: 8], INIT[3454*9 +: 8], INIT[3453*9 +: 8], INIT[3452*9 +: 8], 
          INIT[3451*9 +: 8], INIT[3450*9 +: 8], INIT[3449*9 +: 8], INIT[3448*9 +: 8], 
          INIT[3447*9 +: 8], INIT[3446*9 +: 8], INIT[3445*9 +: 8], INIT[3444*9 +: 8], 
          INIT[3443*9 +: 8], INIT[3442*9 +: 8], INIT[3441*9 +: 8], INIT[3440*9 +: 8], 
          INIT[3439*9 +: 8], INIT[3438*9 +: 8], INIT[3437*9 +: 8], INIT[3436*9 +: 8], 
          INIT[3435*9 +: 8], INIT[3434*9 +: 8], INIT[3433*9 +: 8], INIT[3432*9 +: 8], 
          INIT[3431*9 +: 8], INIT[3430*9 +: 8], INIT[3429*9 +: 8], INIT[3428*9 +: 8], 
          INIT[3427*9 +: 8], INIT[3426*9 +: 8], INIT[3425*9 +: 8], INIT[3424*9 +: 8]}),
.INIT_6C({INIT[3487*9 +: 8], INIT[3486*9 +: 8], INIT[3485*9 +: 8], INIT[3484*9 +: 8], 
          INIT[3483*9 +: 8], INIT[3482*9 +: 8], INIT[3481*9 +: 8], INIT[3480*9 +: 8], 
          INIT[3479*9 +: 8], INIT[3478*9 +: 8], INIT[3477*9 +: 8], INIT[3476*9 +: 8], 
          INIT[3475*9 +: 8], INIT[3474*9 +: 8], INIT[3473*9 +: 8], INIT[3472*9 +: 8], 
          INIT[3471*9 +: 8], INIT[3470*9 +: 8], INIT[3469*9 +: 8], INIT[3468*9 +: 8], 
          INIT[3467*9 +: 8], INIT[3466*9 +: 8], INIT[3465*9 +: 8], INIT[3464*9 +: 8], 
          INIT[3463*9 +: 8], INIT[3462*9 +: 8], INIT[3461*9 +: 8], INIT[3460*9 +: 8], 
          INIT[3459*9 +: 8], INIT[3458*9 +: 8], INIT[3457*9 +: 8], INIT[3456*9 +: 8]}),
.INIT_6D({INIT[3519*9 +: 8], INIT[3518*9 +: 8], INIT[3517*9 +: 8], INIT[3516*9 +: 8], 
          INIT[3515*9 +: 8], INIT[3514*9 +: 8], INIT[3513*9 +: 8], INIT[3512*9 +: 8], 
          INIT[3511*9 +: 8], INIT[3510*9 +: 8], INIT[3509*9 +: 8], INIT[3508*9 +: 8], 
          INIT[3507*9 +: 8], INIT[3506*9 +: 8], INIT[3505*9 +: 8], INIT[3504*9 +: 8], 
          INIT[3503*9 +: 8], INIT[3502*9 +: 8], INIT[3501*9 +: 8], INIT[3500*9 +: 8], 
          INIT[3499*9 +: 8], INIT[3498*9 +: 8], INIT[3497*9 +: 8], INIT[3496*9 +: 8], 
          INIT[3495*9 +: 8], INIT[3494*9 +: 8], INIT[3493*9 +: 8], INIT[3492*9 +: 8], 
          INIT[3491*9 +: 8], INIT[3490*9 +: 8], INIT[3489*9 +: 8], INIT[3488*9 +: 8]}),
.INIT_6E({INIT[3551*9 +: 8], INIT[3550*9 +: 8], INIT[3549*9 +: 8], INIT[3548*9 +: 8], 
          INIT[3547*9 +: 8], INIT[3546*9 +: 8], INIT[3545*9 +: 8], INIT[3544*9 +: 8], 
          INIT[3543*9 +: 8], INIT[3542*9 +: 8], INIT[3541*9 +: 8], INIT[3540*9 +: 8], 
          INIT[3539*9 +: 8], INIT[3538*9 +: 8], INIT[3537*9 +: 8], INIT[3536*9 +: 8], 
          INIT[3535*9 +: 8], INIT[3534*9 +: 8], INIT[3533*9 +: 8], INIT[3532*9 +: 8], 
          INIT[3531*9 +: 8], INIT[3530*9 +: 8], INIT[3529*9 +: 8], INIT[3528*9 +: 8], 
          INIT[3527*9 +: 8], INIT[3526*9 +: 8], INIT[3525*9 +: 8], INIT[3524*9 +: 8], 
          INIT[3523*9 +: 8], INIT[3522*9 +: 8], INIT[3521*9 +: 8], INIT[3520*9 +: 8]}),
.INIT_6F({INIT[3583*9 +: 8], INIT[3582*9 +: 8], INIT[3581*9 +: 8], INIT[3580*9 +: 8], 
          INIT[3579*9 +: 8], INIT[3578*9 +: 8], INIT[3577*9 +: 8], INIT[3576*9 +: 8], 
          INIT[3575*9 +: 8], INIT[3574*9 +: 8], INIT[3573*9 +: 8], INIT[3572*9 +: 8], 
          INIT[3571*9 +: 8], INIT[3570*9 +: 8], INIT[3569*9 +: 8], INIT[3568*9 +: 8], 
          INIT[3567*9 +: 8], INIT[3566*9 +: 8], INIT[3565*9 +: 8], INIT[3564*9 +: 8], 
          INIT[3563*9 +: 8], INIT[3562*9 +: 8], INIT[3561*9 +: 8], INIT[3560*9 +: 8], 
          INIT[3559*9 +: 8], INIT[3558*9 +: 8], INIT[3557*9 +: 8], INIT[3556*9 +: 8], 
          INIT[3555*9 +: 8], INIT[3554*9 +: 8], INIT[3553*9 +: 8], INIT[3552*9 +: 8]}),
.INIT_70({INIT[3615*9 +: 8], INIT[3614*9 +: 8], INIT[3613*9 +: 8], INIT[3612*9 +: 8], 
          INIT[3611*9 +: 8], INIT[3610*9 +: 8], INIT[3609*9 +: 8], INIT[3608*9 +: 8], 
          INIT[3607*9 +: 8], INIT[3606*9 +: 8], INIT[3605*9 +: 8], INIT[3604*9 +: 8], 
          INIT[3603*9 +: 8], INIT[3602*9 +: 8], INIT[3601*9 +: 8], INIT[3600*9 +: 8], 
          INIT[3599*9 +: 8], INIT[3598*9 +: 8], INIT[3597*9 +: 8], INIT[3596*9 +: 8], 
          INIT[3595*9 +: 8], INIT[3594*9 +: 8], INIT[3593*9 +: 8], INIT[3592*9 +: 8], 
          INIT[3591*9 +: 8], INIT[3590*9 +: 8], INIT[3589*9 +: 8], INIT[3588*9 +: 8], 
          INIT[3587*9 +: 8], INIT[3586*9 +: 8], INIT[3585*9 +: 8], INIT[3584*9 +: 8]}),
.INIT_71({INIT[3647*9 +: 8], INIT[3646*9 +: 8], INIT[3645*9 +: 8], INIT[3644*9 +: 8], 
          INIT[3643*9 +: 8], INIT[3642*9 +: 8], INIT[3641*9 +: 8], INIT[3640*9 +: 8], 
          INIT[3639*9 +: 8], INIT[3638*9 +: 8], INIT[3637*9 +: 8], INIT[3636*9 +: 8], 
          INIT[3635*9 +: 8], INIT[3634*9 +: 8], INIT[3633*9 +: 8], INIT[3632*9 +: 8], 
          INIT[3631*9 +: 8], INIT[3630*9 +: 8], INIT[3629*9 +: 8], INIT[3628*9 +: 8], 
          INIT[3627*9 +: 8], INIT[3626*9 +: 8], INIT[3625*9 +: 8], INIT[3624*9 +: 8], 
          INIT[3623*9 +: 8], INIT[3622*9 +: 8], INIT[3621*9 +: 8], INIT[3620*9 +: 8], 
          INIT[3619*9 +: 8], INIT[3618*9 +: 8], INIT[3617*9 +: 8], INIT[3616*9 +: 8]}),
.INIT_72({INIT[3679*9 +: 8], INIT[3678*9 +: 8], INIT[3677*9 +: 8], INIT[3676*9 +: 8], 
          INIT[3675*9 +: 8], INIT[3674*9 +: 8], INIT[3673*9 +: 8], INIT[3672*9 +: 8], 
          INIT[3671*9 +: 8], INIT[3670*9 +: 8], INIT[3669*9 +: 8], INIT[3668*9 +: 8], 
          INIT[3667*9 +: 8], INIT[3666*9 +: 8], INIT[3665*9 +: 8], INIT[3664*9 +: 8], 
          INIT[3663*9 +: 8], INIT[3662*9 +: 8], INIT[3661*9 +: 8], INIT[3660*9 +: 8], 
          INIT[3659*9 +: 8], INIT[3658*9 +: 8], INIT[3657*9 +: 8], INIT[3656*9 +: 8], 
          INIT[3655*9 +: 8], INIT[3654*9 +: 8], INIT[3653*9 +: 8], INIT[3652*9 +: 8], 
          INIT[3651*9 +: 8], INIT[3650*9 +: 8], INIT[3649*9 +: 8], INIT[3648*9 +: 8]}),
.INIT_73({INIT[3711*9 +: 8], INIT[3710*9 +: 8], INIT[3709*9 +: 8], INIT[3708*9 +: 8], 
          INIT[3707*9 +: 8], INIT[3706*9 +: 8], INIT[3705*9 +: 8], INIT[3704*9 +: 8], 
          INIT[3703*9 +: 8], INIT[3702*9 +: 8], INIT[3701*9 +: 8], INIT[3700*9 +: 8], 
          INIT[3699*9 +: 8], INIT[3698*9 +: 8], INIT[3697*9 +: 8], INIT[3696*9 +: 8], 
          INIT[3695*9 +: 8], INIT[3694*9 +: 8], INIT[3693*9 +: 8], INIT[3692*9 +: 8], 
          INIT[3691*9 +: 8], INIT[3690*9 +: 8], INIT[3689*9 +: 8], INIT[3688*9 +: 8], 
          INIT[3687*9 +: 8], INIT[3686*9 +: 8], INIT[3685*9 +: 8], INIT[3684*9 +: 8], 
          INIT[3683*9 +: 8], INIT[3682*9 +: 8], INIT[3681*9 +: 8], INIT[3680*9 +: 8]}),
.INIT_74({INIT[3743*9 +: 8], INIT[3742*9 +: 8], INIT[3741*9 +: 8], INIT[3740*9 +: 8], 
          INIT[3739*9 +: 8], INIT[3738*9 +: 8], INIT[3737*9 +: 8], INIT[3736*9 +: 8], 
          INIT[3735*9 +: 8], INIT[3734*9 +: 8], INIT[3733*9 +: 8], INIT[3732*9 +: 8], 
          INIT[3731*9 +: 8], INIT[3730*9 +: 8], INIT[3729*9 +: 8], INIT[3728*9 +: 8], 
          INIT[3727*9 +: 8], INIT[3726*9 +: 8], INIT[3725*9 +: 8], INIT[3724*9 +: 8], 
          INIT[3723*9 +: 8], INIT[3722*9 +: 8], INIT[3721*9 +: 8], INIT[3720*9 +: 8], 
          INIT[3719*9 +: 8], INIT[3718*9 +: 8], INIT[3717*9 +: 8], INIT[3716*9 +: 8], 
          INIT[3715*9 +: 8], INIT[3714*9 +: 8], INIT[3713*9 +: 8], INIT[3712*9 +: 8]}),
.INIT_75({INIT[3775*9 +: 8], INIT[3774*9 +: 8], INIT[3773*9 +: 8], INIT[3772*9 +: 8], 
          INIT[3771*9 +: 8], INIT[3770*9 +: 8], INIT[3769*9 +: 8], INIT[3768*9 +: 8], 
          INIT[3767*9 +: 8], INIT[3766*9 +: 8], INIT[3765*9 +: 8], INIT[3764*9 +: 8], 
          INIT[3763*9 +: 8], INIT[3762*9 +: 8], INIT[3761*9 +: 8], INIT[3760*9 +: 8], 
          INIT[3759*9 +: 8], INIT[3758*9 +: 8], INIT[3757*9 +: 8], INIT[3756*9 +: 8], 
          INIT[3755*9 +: 8], INIT[3754*9 +: 8], INIT[3753*9 +: 8], INIT[3752*9 +: 8], 
          INIT[3751*9 +: 8], INIT[3750*9 +: 8], INIT[3749*9 +: 8], INIT[3748*9 +: 8], 
          INIT[3747*9 +: 8], INIT[3746*9 +: 8], INIT[3745*9 +: 8], INIT[3744*9 +: 8]}),
.INIT_76({INIT[3807*9 +: 8], INIT[3806*9 +: 8], INIT[3805*9 +: 8], INIT[3804*9 +: 8], 
          INIT[3803*9 +: 8], INIT[3802*9 +: 8], INIT[3801*9 +: 8], INIT[3800*9 +: 8], 
          INIT[3799*9 +: 8], INIT[3798*9 +: 8], INIT[3797*9 +: 8], INIT[3796*9 +: 8], 
          INIT[3795*9 +: 8], INIT[3794*9 +: 8], INIT[3793*9 +: 8], INIT[3792*9 +: 8], 
          INIT[3791*9 +: 8], INIT[3790*9 +: 8], INIT[3789*9 +: 8], INIT[3788*9 +: 8], 
          INIT[3787*9 +: 8], INIT[3786*9 +: 8], INIT[3785*9 +: 8], INIT[3784*9 +: 8], 
          INIT[3783*9 +: 8], INIT[3782*9 +: 8], INIT[3781*9 +: 8], INIT[3780*9 +: 8], 
          INIT[3779*9 +: 8], INIT[3778*9 +: 8], INIT[3777*9 +: 8], INIT[3776*9 +: 8]}),
.INIT_77({INIT[3839*9 +: 8], INIT[3838*9 +: 8], INIT[3837*9 +: 8], INIT[3836*9 +: 8], 
          INIT[3835*9 +: 8], INIT[3834*9 +: 8], INIT[3833*9 +: 8], INIT[3832*9 +: 8], 
          INIT[3831*9 +: 8], INIT[3830*9 +: 8], INIT[3829*9 +: 8], INIT[3828*9 +: 8], 
          INIT[3827*9 +: 8], INIT[3826*9 +: 8], INIT[3825*9 +: 8], INIT[3824*9 +: 8], 
          INIT[3823*9 +: 8], INIT[3822*9 +: 8], INIT[3821*9 +: 8], INIT[3820*9 +: 8], 
          INIT[3819*9 +: 8], INIT[3818*9 +: 8], INIT[3817*9 +: 8], INIT[3816*9 +: 8], 
          INIT[3815*9 +: 8], INIT[3814*9 +: 8], INIT[3813*9 +: 8], INIT[3812*9 +: 8], 
          INIT[3811*9 +: 8], INIT[3810*9 +: 8], INIT[3809*9 +: 8], INIT[3808*9 +: 8]}),
.INIT_78({INIT[3871*9 +: 8], INIT[3870*9 +: 8], INIT[3869*9 +: 8], INIT[3868*9 +: 8], 
          INIT[3867*9 +: 8], INIT[3866*9 +: 8], INIT[3865*9 +: 8], INIT[3864*9 +: 8], 
          INIT[3863*9 +: 8], INIT[3862*9 +: 8], INIT[3861*9 +: 8], INIT[3860*9 +: 8], 
          INIT[3859*9 +: 8], INIT[3858*9 +: 8], INIT[3857*9 +: 8], INIT[3856*9 +: 8], 
          INIT[3855*9 +: 8], INIT[3854*9 +: 8], INIT[3853*9 +: 8], INIT[3852*9 +: 8], 
          INIT[3851*9 +: 8], INIT[3850*9 +: 8], INIT[3849*9 +: 8], INIT[3848*9 +: 8], 
          INIT[3847*9 +: 8], INIT[3846*9 +: 8], INIT[3845*9 +: 8], INIT[3844*9 +: 8], 
          INIT[3843*9 +: 8], INIT[3842*9 +: 8], INIT[3841*9 +: 8], INIT[3840*9 +: 8]}),
.INIT_79({INIT[3903*9 +: 8], INIT[3902*9 +: 8], INIT[3901*9 +: 8], INIT[3900*9 +: 8], 
          INIT[3899*9 +: 8], INIT[3898*9 +: 8], INIT[3897*9 +: 8], INIT[3896*9 +: 8], 
          INIT[3895*9 +: 8], INIT[3894*9 +: 8], INIT[3893*9 +: 8], INIT[3892*9 +: 8], 
          INIT[3891*9 +: 8], INIT[3890*9 +: 8], INIT[3889*9 +: 8], INIT[3888*9 +: 8], 
          INIT[3887*9 +: 8], INIT[3886*9 +: 8], INIT[3885*9 +: 8], INIT[3884*9 +: 8], 
          INIT[3883*9 +: 8], INIT[3882*9 +: 8], INIT[3881*9 +: 8], INIT[3880*9 +: 8], 
          INIT[3879*9 +: 8], INIT[3878*9 +: 8], INIT[3877*9 +: 8], INIT[3876*9 +: 8], 
          INIT[3875*9 +: 8], INIT[3874*9 +: 8], INIT[3873*9 +: 8], INIT[3872*9 +: 8]}),
.INIT_7A({INIT[3935*9 +: 8], INIT[3934*9 +: 8], INIT[3933*9 +: 8], INIT[3932*9 +: 8], 
          INIT[3931*9 +: 8], INIT[3930*9 +: 8], INIT[3929*9 +: 8], INIT[3928*9 +: 8], 
          INIT[3927*9 +: 8], INIT[3926*9 +: 8], INIT[3925*9 +: 8], INIT[3924*9 +: 8], 
          INIT[3923*9 +: 8], INIT[3922*9 +: 8], INIT[3921*9 +: 8], INIT[3920*9 +: 8], 
          INIT[3919*9 +: 8], INIT[3918*9 +: 8], INIT[3917*9 +: 8], INIT[3916*9 +: 8], 
          INIT[3915*9 +: 8], INIT[3914*9 +: 8], INIT[3913*9 +: 8], INIT[3912*9 +: 8], 
          INIT[3911*9 +: 8], INIT[3910*9 +: 8], INIT[3909*9 +: 8], INIT[3908*9 +: 8], 
          INIT[3907*9 +: 8], INIT[3906*9 +: 8], INIT[3905*9 +: 8], INIT[3904*9 +: 8]}),
.INIT_7B({INIT[3967*9 +: 8], INIT[3966*9 +: 8], INIT[3965*9 +: 8], INIT[3964*9 +: 8], 
          INIT[3963*9 +: 8], INIT[3962*9 +: 8], INIT[3961*9 +: 8], INIT[3960*9 +: 8], 
          INIT[3959*9 +: 8], INIT[3958*9 +: 8], INIT[3957*9 +: 8], INIT[3956*9 +: 8], 
          INIT[3955*9 +: 8], INIT[3954*9 +: 8], INIT[3953*9 +: 8], INIT[3952*9 +: 8], 
          INIT[3951*9 +: 8], INIT[3950*9 +: 8], INIT[3949*9 +: 8], INIT[3948*9 +: 8], 
          INIT[3947*9 +: 8], INIT[3946*9 +: 8], INIT[3945*9 +: 8], INIT[3944*9 +: 8], 
          INIT[3943*9 +: 8], INIT[3942*9 +: 8], INIT[3941*9 +: 8], INIT[3940*9 +: 8], 
          INIT[3939*9 +: 8], INIT[3938*9 +: 8], INIT[3937*9 +: 8], INIT[3936*9 +: 8]}),
.INIT_7C({INIT[3999*9 +: 8], INIT[3998*9 +: 8], INIT[3997*9 +: 8], INIT[3996*9 +: 8], 
          INIT[3995*9 +: 8], INIT[3994*9 +: 8], INIT[3993*9 +: 8], INIT[3992*9 +: 8], 
          INIT[3991*9 +: 8], INIT[3990*9 +: 8], INIT[3989*9 +: 8], INIT[3988*9 +: 8], 
          INIT[3987*9 +: 8], INIT[3986*9 +: 8], INIT[3985*9 +: 8], INIT[3984*9 +: 8], 
          INIT[3983*9 +: 8], INIT[3982*9 +: 8], INIT[3981*9 +: 8], INIT[3980*9 +: 8], 
          INIT[3979*9 +: 8], INIT[3978*9 +: 8], INIT[3977*9 +: 8], INIT[3976*9 +: 8], 
          INIT[3975*9 +: 8], INIT[3974*9 +: 8], INIT[3973*9 +: 8], INIT[3972*9 +: 8], 
          INIT[3971*9 +: 8], INIT[3970*9 +: 8], INIT[3969*9 +: 8], INIT[3968*9 +: 8]}),
.INIT_7D({INIT[4031*9 +: 8], INIT[4030*9 +: 8], INIT[4029*9 +: 8], INIT[4028*9 +: 8], 
          INIT[4027*9 +: 8], INIT[4026*9 +: 8], INIT[4025*9 +: 8], INIT[4024*9 +: 8], 
          INIT[4023*9 +: 8], INIT[4022*9 +: 8], INIT[4021*9 +: 8], INIT[4020*9 +: 8], 
          INIT[4019*9 +: 8], INIT[4018*9 +: 8], INIT[4017*9 +: 8], INIT[4016*9 +: 8], 
          INIT[4015*9 +: 8], INIT[4014*9 +: 8], INIT[4013*9 +: 8], INIT[4012*9 +: 8], 
          INIT[4011*9 +: 8], INIT[4010*9 +: 8], INIT[4009*9 +: 8], INIT[4008*9 +: 8], 
          INIT[4007*9 +: 8], INIT[4006*9 +: 8], INIT[4005*9 +: 8], INIT[4004*9 +: 8], 
          INIT[4003*9 +: 8], INIT[4002*9 +: 8], INIT[4001*9 +: 8], INIT[4000*9 +: 8]}),
.INIT_7E({INIT[4063*9 +: 8], INIT[4062*9 +: 8], INIT[4061*9 +: 8], INIT[4060*9 +: 8], 
          INIT[4059*9 +: 8], INIT[4058*9 +: 8], INIT[4057*9 +: 8], INIT[4056*9 +: 8], 
          INIT[4055*9 +: 8], INIT[4054*9 +: 8], INIT[4053*9 +: 8], INIT[4052*9 +: 8], 
          INIT[4051*9 +: 8], INIT[4050*9 +: 8], INIT[4049*9 +: 8], INIT[4048*9 +: 8], 
          INIT[4047*9 +: 8], INIT[4046*9 +: 8], INIT[4045*9 +: 8], INIT[4044*9 +: 8], 
          INIT[4043*9 +: 8], INIT[4042*9 +: 8], INIT[4041*9 +: 8], INIT[4040*9 +: 8], 
          INIT[4039*9 +: 8], INIT[4038*9 +: 8], INIT[4037*9 +: 8], INIT[4036*9 +: 8], 
          INIT[4035*9 +: 8], INIT[4034*9 +: 8], INIT[4033*9 +: 8], INIT[4032*9 +: 8]}),
.INIT_7F({INIT[4095*9 +: 8], INIT[4094*9 +: 8], INIT[4093*9 +: 8], INIT[4092*9 +: 8], 
          INIT[4091*9 +: 8], INIT[4090*9 +: 8], INIT[4089*9 +: 8], INIT[4088*9 +: 8], 
          INIT[4087*9 +: 8], INIT[4086*9 +: 8], INIT[4085*9 +: 8], INIT[4084*9 +: 8], 
          INIT[4083*9 +: 8], INIT[4082*9 +: 8], INIT[4081*9 +: 8], INIT[4080*9 +: 8], 
          INIT[4079*9 +: 8], INIT[4078*9 +: 8], INIT[4077*9 +: 8], INIT[4076*9 +: 8], 
          INIT[4075*9 +: 8], INIT[4074*9 +: 8], INIT[4073*9 +: 8], INIT[4072*9 +: 8], 
          INIT[4071*9 +: 8], INIT[4070*9 +: 8], INIT[4069*9 +: 8], INIT[4068*9 +: 8], 
          INIT[4067*9 +: 8], INIT[4066*9 +: 8], INIT[4065*9 +: 8], INIT[4064*9 +: 8]}),
