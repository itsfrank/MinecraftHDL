.INIT_00(INIT[  0*256 +: 256]),
.INIT_01(INIT[  1*256 +: 256]),
.INIT_02(INIT[  2*256 +: 256]),
.INIT_03(INIT[  3*256 +: 256]),
.INIT_04(INIT[  4*256 +: 256]),
.INIT_05(INIT[  5*256 +: 256]),
.INIT_06(INIT[  6*256 +: 256]),
.INIT_07(INIT[  7*256 +: 256]),
.INIT_08(INIT[  8*256 +: 256]),
.INIT_09(INIT[  9*256 +: 256]),
.INIT_0A(INIT[ 10*256 +: 256]),
.INIT_0B(INIT[ 11*256 +: 256]),
.INIT_0C(INIT[ 12*256 +: 256]),
.INIT_0D(INIT[ 13*256 +: 256]),
.INIT_0E(INIT[ 14*256 +: 256]),
.INIT_0F(INIT[ 15*256 +: 256]),
.INIT_10(INIT[ 16*256 +: 256]),
.INIT_11(INIT[ 17*256 +: 256]),
.INIT_12(INIT[ 18*256 +: 256]),
.INIT_13(INIT[ 19*256 +: 256]),
.INIT_14(INIT[ 20*256 +: 256]),
.INIT_15(INIT[ 21*256 +: 256]),
.INIT_16(INIT[ 22*256 +: 256]),
.INIT_17(INIT[ 23*256 +: 256]),
.INIT_18(INIT[ 24*256 +: 256]),
.INIT_19(INIT[ 25*256 +: 256]),
.INIT_1A(INIT[ 26*256 +: 256]),
.INIT_1B(INIT[ 27*256 +: 256]),
.INIT_1C(INIT[ 28*256 +: 256]),
.INIT_1D(INIT[ 29*256 +: 256]),
.INIT_1E(INIT[ 30*256 +: 256]),
.INIT_1F(INIT[ 31*256 +: 256]),
.INIT_20(INIT[ 32*256 +: 256]),
.INIT_21(INIT[ 33*256 +: 256]),
.INIT_22(INIT[ 34*256 +: 256]),
.INIT_23(INIT[ 35*256 +: 256]),
.INIT_24(INIT[ 36*256 +: 256]),
.INIT_25(INIT[ 37*256 +: 256]),
.INIT_26(INIT[ 38*256 +: 256]),
.INIT_27(INIT[ 39*256 +: 256]),
.INIT_28(INIT[ 40*256 +: 256]),
.INIT_29(INIT[ 41*256 +: 256]),
.INIT_2A(INIT[ 42*256 +: 256]),
.INIT_2B(INIT[ 43*256 +: 256]),
.INIT_2C(INIT[ 44*256 +: 256]),
.INIT_2D(INIT[ 45*256 +: 256]),
.INIT_2E(INIT[ 46*256 +: 256]),
.INIT_2F(INIT[ 47*256 +: 256]),
.INIT_30(INIT[ 48*256 +: 256]),
.INIT_31(INIT[ 49*256 +: 256]),
.INIT_32(INIT[ 50*256 +: 256]),
.INIT_33(INIT[ 51*256 +: 256]),
.INIT_34(INIT[ 52*256 +: 256]),
.INIT_35(INIT[ 53*256 +: 256]),
.INIT_36(INIT[ 54*256 +: 256]),
.INIT_37(INIT[ 55*256 +: 256]),
.INIT_38(INIT[ 56*256 +: 256]),
.INIT_39(INIT[ 57*256 +: 256]),
.INIT_3A(INIT[ 58*256 +: 256]),
.INIT_3B(INIT[ 59*256 +: 256]),
.INIT_3C(INIT[ 60*256 +: 256]),
.INIT_3D(INIT[ 61*256 +: 256]),
.INIT_3E(INIT[ 62*256 +: 256]),
.INIT_3F(INIT[ 63*256 +: 256]),
.INIT_40(INIT[ 64*256 +: 256]),
.INIT_41(INIT[ 65*256 +: 256]),
.INIT_42(INIT[ 66*256 +: 256]),
.INIT_43(INIT[ 67*256 +: 256]),
.INIT_44(INIT[ 68*256 +: 256]),
.INIT_45(INIT[ 69*256 +: 256]),
.INIT_46(INIT[ 70*256 +: 256]),
.INIT_47(INIT[ 71*256 +: 256]),
.INIT_48(INIT[ 72*256 +: 256]),
.INIT_49(INIT[ 73*256 +: 256]),
.INIT_4A(INIT[ 74*256 +: 256]),
.INIT_4B(INIT[ 75*256 +: 256]),
.INIT_4C(INIT[ 76*256 +: 256]),
.INIT_4D(INIT[ 77*256 +: 256]),
.INIT_4E(INIT[ 78*256 +: 256]),
.INIT_4F(INIT[ 79*256 +: 256]),
.INIT_50(INIT[ 80*256 +: 256]),
.INIT_51(INIT[ 81*256 +: 256]),
.INIT_52(INIT[ 82*256 +: 256]),
.INIT_53(INIT[ 83*256 +: 256]),
.INIT_54(INIT[ 84*256 +: 256]),
.INIT_55(INIT[ 85*256 +: 256]),
.INIT_56(INIT[ 86*256 +: 256]),
.INIT_57(INIT[ 87*256 +: 256]),
.INIT_58(INIT[ 88*256 +: 256]),
.INIT_59(INIT[ 89*256 +: 256]),
.INIT_5A(INIT[ 90*256 +: 256]),
.INIT_5B(INIT[ 91*256 +: 256]),
.INIT_5C(INIT[ 92*256 +: 256]),
.INIT_5D(INIT[ 93*256 +: 256]),
.INIT_5E(INIT[ 94*256 +: 256]),
.INIT_5F(INIT[ 95*256 +: 256]),
.INIT_60(INIT[ 96*256 +: 256]),
.INIT_61(INIT[ 97*256 +: 256]),
.INIT_62(INIT[ 98*256 +: 256]),
.INIT_63(INIT[ 99*256 +: 256]),
.INIT_64(INIT[100*256 +: 256]),
.INIT_65(INIT[101*256 +: 256]),
.INIT_66(INIT[102*256 +: 256]),
.INIT_67(INIT[103*256 +: 256]),
.INIT_68(INIT[104*256 +: 256]),
.INIT_69(INIT[105*256 +: 256]),
.INIT_6A(INIT[106*256 +: 256]),
.INIT_6B(INIT[107*256 +: 256]),
.INIT_6C(INIT[108*256 +: 256]),
.INIT_6D(INIT[109*256 +: 256]),
.INIT_6E(INIT[110*256 +: 256]),
.INIT_6F(INIT[111*256 +: 256]),
.INIT_70(INIT[112*256 +: 256]),
.INIT_71(INIT[113*256 +: 256]),
.INIT_72(INIT[114*256 +: 256]),
.INIT_73(INIT[115*256 +: 256]),
.INIT_74(INIT[116*256 +: 256]),
.INIT_75(INIT[117*256 +: 256]),
.INIT_76(INIT[118*256 +: 256]),
.INIT_77(INIT[119*256 +: 256]),
.INIT_78(INIT[120*256 +: 256]),
.INIT_79(INIT[121*256 +: 256]),
.INIT_7A(INIT[122*256 +: 256]),
.INIT_7B(INIT[123*256 +: 256]),
.INIT_7C(INIT[124*256 +: 256]),
.INIT_7D(INIT[125*256 +: 256]),
.INIT_7E(INIT[126*256 +: 256]),
.INIT_7F(INIT[127*256 +: 256]),
