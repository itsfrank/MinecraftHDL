module OR(a, b, c, out);
input a, b, c;
output out;
OR G1(out, a, b, c);
endmodule