module testAND(input a, input b, output c);
AND G1(c, a, b);
endmodule

