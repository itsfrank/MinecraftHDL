localparam [255:0] INIT_0 = {
  INIT[3615], INIT[3103], INIT[2591], INIT[2079], INIT[1567], INIT[1055], INIT[ 543], INIT[  31],
  INIT[3614], INIT[3102], INIT[2590], INIT[2078], INIT[1566], INIT[1054], INIT[ 542], INIT[  30],
  INIT[3613], INIT[3101], INIT[2589], INIT[2077], INIT[1565], INIT[1053], INIT[ 541], INIT[  29],
  INIT[3612], INIT[3100], INIT[2588], INIT[2076], INIT[1564], INIT[1052], INIT[ 540], INIT[  28],
  INIT[3611], INIT[3099], INIT[2587], INIT[2075], INIT[1563], INIT[1051], INIT[ 539], INIT[  27],
  INIT[3610], INIT[3098], INIT[2586], INIT[2074], INIT[1562], INIT[1050], INIT[ 538], INIT[  26],
  INIT[3609], INIT[3097], INIT[2585], INIT[2073], INIT[1561], INIT[1049], INIT[ 537], INIT[  25],
  INIT[3608], INIT[3096], INIT[2584], INIT[2072], INIT[1560], INIT[1048], INIT[ 536], INIT[  24],
  INIT[3607], INIT[3095], INIT[2583], INIT[2071], INIT[1559], INIT[1047], INIT[ 535], INIT[  23],
  INIT[3606], INIT[3094], INIT[2582], INIT[2070], INIT[1558], INIT[1046], INIT[ 534], INIT[  22],
  INIT[3605], INIT[3093], INIT[2581], INIT[2069], INIT[1557], INIT[1045], INIT[ 533], INIT[  21],
  INIT[3604], INIT[3092], INIT[2580], INIT[2068], INIT[1556], INIT[1044], INIT[ 532], INIT[  20],
  INIT[3603], INIT[3091], INIT[2579], INIT[2067], INIT[1555], INIT[1043], INIT[ 531], INIT[  19],
  INIT[3602], INIT[3090], INIT[2578], INIT[2066], INIT[1554], INIT[1042], INIT[ 530], INIT[  18],
  INIT[3601], INIT[3089], INIT[2577], INIT[2065], INIT[1553], INIT[1041], INIT[ 529], INIT[  17],
  INIT[3600], INIT[3088], INIT[2576], INIT[2064], INIT[1552], INIT[1040], INIT[ 528], INIT[  16],
  INIT[3599], INIT[3087], INIT[2575], INIT[2063], INIT[1551], INIT[1039], INIT[ 527], INIT[  15],
  INIT[3598], INIT[3086], INIT[2574], INIT[2062], INIT[1550], INIT[1038], INIT[ 526], INIT[  14],
  INIT[3597], INIT[3085], INIT[2573], INIT[2061], INIT[1549], INIT[1037], INIT[ 525], INIT[  13],
  INIT[3596], INIT[3084], INIT[2572], INIT[2060], INIT[1548], INIT[1036], INIT[ 524], INIT[  12],
  INIT[3595], INIT[3083], INIT[2571], INIT[2059], INIT[1547], INIT[1035], INIT[ 523], INIT[  11],
  INIT[3594], INIT[3082], INIT[2570], INIT[2058], INIT[1546], INIT[1034], INIT[ 522], INIT[  10],
  INIT[3593], INIT[3081], INIT[2569], INIT[2057], INIT[1545], INIT[1033], INIT[ 521], INIT[   9],
  INIT[3592], INIT[3080], INIT[2568], INIT[2056], INIT[1544], INIT[1032], INIT[ 520], INIT[   8],
  INIT[3591], INIT[3079], INIT[2567], INIT[2055], INIT[1543], INIT[1031], INIT[ 519], INIT[   7],
  INIT[3590], INIT[3078], INIT[2566], INIT[2054], INIT[1542], INIT[1030], INIT[ 518], INIT[   6],
  INIT[3589], INIT[3077], INIT[2565], INIT[2053], INIT[1541], INIT[1029], INIT[ 517], INIT[   5],
  INIT[3588], INIT[3076], INIT[2564], INIT[2052], INIT[1540], INIT[1028], INIT[ 516], INIT[   4],
  INIT[3587], INIT[3075], INIT[2563], INIT[2051], INIT[1539], INIT[1027], INIT[ 515], INIT[   3],
  INIT[3586], INIT[3074], INIT[2562], INIT[2050], INIT[1538], INIT[1026], INIT[ 514], INIT[   2],
  INIT[3585], INIT[3073], INIT[2561], INIT[2049], INIT[1537], INIT[1025], INIT[ 513], INIT[   1],
  INIT[3584], INIT[3072], INIT[2560], INIT[2048], INIT[1536], INIT[1024], INIT[ 512], INIT[   0]
};
localparam [255:0] INIT_1 = {
  INIT[3647], INIT[3135], INIT[2623], INIT[2111], INIT[1599], INIT[1087], INIT[ 575], INIT[  63],
  INIT[3646], INIT[3134], INIT[2622], INIT[2110], INIT[1598], INIT[1086], INIT[ 574], INIT[  62],
  INIT[3645], INIT[3133], INIT[2621], INIT[2109], INIT[1597], INIT[1085], INIT[ 573], INIT[  61],
  INIT[3644], INIT[3132], INIT[2620], INIT[2108], INIT[1596], INIT[1084], INIT[ 572], INIT[  60],
  INIT[3643], INIT[3131], INIT[2619], INIT[2107], INIT[1595], INIT[1083], INIT[ 571], INIT[  59],
  INIT[3642], INIT[3130], INIT[2618], INIT[2106], INIT[1594], INIT[1082], INIT[ 570], INIT[  58],
  INIT[3641], INIT[3129], INIT[2617], INIT[2105], INIT[1593], INIT[1081], INIT[ 569], INIT[  57],
  INIT[3640], INIT[3128], INIT[2616], INIT[2104], INIT[1592], INIT[1080], INIT[ 568], INIT[  56],
  INIT[3639], INIT[3127], INIT[2615], INIT[2103], INIT[1591], INIT[1079], INIT[ 567], INIT[  55],
  INIT[3638], INIT[3126], INIT[2614], INIT[2102], INIT[1590], INIT[1078], INIT[ 566], INIT[  54],
  INIT[3637], INIT[3125], INIT[2613], INIT[2101], INIT[1589], INIT[1077], INIT[ 565], INIT[  53],
  INIT[3636], INIT[3124], INIT[2612], INIT[2100], INIT[1588], INIT[1076], INIT[ 564], INIT[  52],
  INIT[3635], INIT[3123], INIT[2611], INIT[2099], INIT[1587], INIT[1075], INIT[ 563], INIT[  51],
  INIT[3634], INIT[3122], INIT[2610], INIT[2098], INIT[1586], INIT[1074], INIT[ 562], INIT[  50],
  INIT[3633], INIT[3121], INIT[2609], INIT[2097], INIT[1585], INIT[1073], INIT[ 561], INIT[  49],
  INIT[3632], INIT[3120], INIT[2608], INIT[2096], INIT[1584], INIT[1072], INIT[ 560], INIT[  48],
  INIT[3631], INIT[3119], INIT[2607], INIT[2095], INIT[1583], INIT[1071], INIT[ 559], INIT[  47],
  INIT[3630], INIT[3118], INIT[2606], INIT[2094], INIT[1582], INIT[1070], INIT[ 558], INIT[  46],
  INIT[3629], INIT[3117], INIT[2605], INIT[2093], INIT[1581], INIT[1069], INIT[ 557], INIT[  45],
  INIT[3628], INIT[3116], INIT[2604], INIT[2092], INIT[1580], INIT[1068], INIT[ 556], INIT[  44],
  INIT[3627], INIT[3115], INIT[2603], INIT[2091], INIT[1579], INIT[1067], INIT[ 555], INIT[  43],
  INIT[3626], INIT[3114], INIT[2602], INIT[2090], INIT[1578], INIT[1066], INIT[ 554], INIT[  42],
  INIT[3625], INIT[3113], INIT[2601], INIT[2089], INIT[1577], INIT[1065], INIT[ 553], INIT[  41],
  INIT[3624], INIT[3112], INIT[2600], INIT[2088], INIT[1576], INIT[1064], INIT[ 552], INIT[  40],
  INIT[3623], INIT[3111], INIT[2599], INIT[2087], INIT[1575], INIT[1063], INIT[ 551], INIT[  39],
  INIT[3622], INIT[3110], INIT[2598], INIT[2086], INIT[1574], INIT[1062], INIT[ 550], INIT[  38],
  INIT[3621], INIT[3109], INIT[2597], INIT[2085], INIT[1573], INIT[1061], INIT[ 549], INIT[  37],
  INIT[3620], INIT[3108], INIT[2596], INIT[2084], INIT[1572], INIT[1060], INIT[ 548], INIT[  36],
  INIT[3619], INIT[3107], INIT[2595], INIT[2083], INIT[1571], INIT[1059], INIT[ 547], INIT[  35],
  INIT[3618], INIT[3106], INIT[2594], INIT[2082], INIT[1570], INIT[1058], INIT[ 546], INIT[  34],
  INIT[3617], INIT[3105], INIT[2593], INIT[2081], INIT[1569], INIT[1057], INIT[ 545], INIT[  33],
  INIT[3616], INIT[3104], INIT[2592], INIT[2080], INIT[1568], INIT[1056], INIT[ 544], INIT[  32]
};
localparam [255:0] INIT_2 = {
  INIT[3679], INIT[3167], INIT[2655], INIT[2143], INIT[1631], INIT[1119], INIT[ 607], INIT[  95],
  INIT[3678], INIT[3166], INIT[2654], INIT[2142], INIT[1630], INIT[1118], INIT[ 606], INIT[  94],
  INIT[3677], INIT[3165], INIT[2653], INIT[2141], INIT[1629], INIT[1117], INIT[ 605], INIT[  93],
  INIT[3676], INIT[3164], INIT[2652], INIT[2140], INIT[1628], INIT[1116], INIT[ 604], INIT[  92],
  INIT[3675], INIT[3163], INIT[2651], INIT[2139], INIT[1627], INIT[1115], INIT[ 603], INIT[  91],
  INIT[3674], INIT[3162], INIT[2650], INIT[2138], INIT[1626], INIT[1114], INIT[ 602], INIT[  90],
  INIT[3673], INIT[3161], INIT[2649], INIT[2137], INIT[1625], INIT[1113], INIT[ 601], INIT[  89],
  INIT[3672], INIT[3160], INIT[2648], INIT[2136], INIT[1624], INIT[1112], INIT[ 600], INIT[  88],
  INIT[3671], INIT[3159], INIT[2647], INIT[2135], INIT[1623], INIT[1111], INIT[ 599], INIT[  87],
  INIT[3670], INIT[3158], INIT[2646], INIT[2134], INIT[1622], INIT[1110], INIT[ 598], INIT[  86],
  INIT[3669], INIT[3157], INIT[2645], INIT[2133], INIT[1621], INIT[1109], INIT[ 597], INIT[  85],
  INIT[3668], INIT[3156], INIT[2644], INIT[2132], INIT[1620], INIT[1108], INIT[ 596], INIT[  84],
  INIT[3667], INIT[3155], INIT[2643], INIT[2131], INIT[1619], INIT[1107], INIT[ 595], INIT[  83],
  INIT[3666], INIT[3154], INIT[2642], INIT[2130], INIT[1618], INIT[1106], INIT[ 594], INIT[  82],
  INIT[3665], INIT[3153], INIT[2641], INIT[2129], INIT[1617], INIT[1105], INIT[ 593], INIT[  81],
  INIT[3664], INIT[3152], INIT[2640], INIT[2128], INIT[1616], INIT[1104], INIT[ 592], INIT[  80],
  INIT[3663], INIT[3151], INIT[2639], INIT[2127], INIT[1615], INIT[1103], INIT[ 591], INIT[  79],
  INIT[3662], INIT[3150], INIT[2638], INIT[2126], INIT[1614], INIT[1102], INIT[ 590], INIT[  78],
  INIT[3661], INIT[3149], INIT[2637], INIT[2125], INIT[1613], INIT[1101], INIT[ 589], INIT[  77],
  INIT[3660], INIT[3148], INIT[2636], INIT[2124], INIT[1612], INIT[1100], INIT[ 588], INIT[  76],
  INIT[3659], INIT[3147], INIT[2635], INIT[2123], INIT[1611], INIT[1099], INIT[ 587], INIT[  75],
  INIT[3658], INIT[3146], INIT[2634], INIT[2122], INIT[1610], INIT[1098], INIT[ 586], INIT[  74],
  INIT[3657], INIT[3145], INIT[2633], INIT[2121], INIT[1609], INIT[1097], INIT[ 585], INIT[  73],
  INIT[3656], INIT[3144], INIT[2632], INIT[2120], INIT[1608], INIT[1096], INIT[ 584], INIT[  72],
  INIT[3655], INIT[3143], INIT[2631], INIT[2119], INIT[1607], INIT[1095], INIT[ 583], INIT[  71],
  INIT[3654], INIT[3142], INIT[2630], INIT[2118], INIT[1606], INIT[1094], INIT[ 582], INIT[  70],
  INIT[3653], INIT[3141], INIT[2629], INIT[2117], INIT[1605], INIT[1093], INIT[ 581], INIT[  69],
  INIT[3652], INIT[3140], INIT[2628], INIT[2116], INIT[1604], INIT[1092], INIT[ 580], INIT[  68],
  INIT[3651], INIT[3139], INIT[2627], INIT[2115], INIT[1603], INIT[1091], INIT[ 579], INIT[  67],
  INIT[3650], INIT[3138], INIT[2626], INIT[2114], INIT[1602], INIT[1090], INIT[ 578], INIT[  66],
  INIT[3649], INIT[3137], INIT[2625], INIT[2113], INIT[1601], INIT[1089], INIT[ 577], INIT[  65],
  INIT[3648], INIT[3136], INIT[2624], INIT[2112], INIT[1600], INIT[1088], INIT[ 576], INIT[  64]
};
localparam [255:0] INIT_3 = {
  INIT[3711], INIT[3199], INIT[2687], INIT[2175], INIT[1663], INIT[1151], INIT[ 639], INIT[ 127],
  INIT[3710], INIT[3198], INIT[2686], INIT[2174], INIT[1662], INIT[1150], INIT[ 638], INIT[ 126],
  INIT[3709], INIT[3197], INIT[2685], INIT[2173], INIT[1661], INIT[1149], INIT[ 637], INIT[ 125],
  INIT[3708], INIT[3196], INIT[2684], INIT[2172], INIT[1660], INIT[1148], INIT[ 636], INIT[ 124],
  INIT[3707], INIT[3195], INIT[2683], INIT[2171], INIT[1659], INIT[1147], INIT[ 635], INIT[ 123],
  INIT[3706], INIT[3194], INIT[2682], INIT[2170], INIT[1658], INIT[1146], INIT[ 634], INIT[ 122],
  INIT[3705], INIT[3193], INIT[2681], INIT[2169], INIT[1657], INIT[1145], INIT[ 633], INIT[ 121],
  INIT[3704], INIT[3192], INIT[2680], INIT[2168], INIT[1656], INIT[1144], INIT[ 632], INIT[ 120],
  INIT[3703], INIT[3191], INIT[2679], INIT[2167], INIT[1655], INIT[1143], INIT[ 631], INIT[ 119],
  INIT[3702], INIT[3190], INIT[2678], INIT[2166], INIT[1654], INIT[1142], INIT[ 630], INIT[ 118],
  INIT[3701], INIT[3189], INIT[2677], INIT[2165], INIT[1653], INIT[1141], INIT[ 629], INIT[ 117],
  INIT[3700], INIT[3188], INIT[2676], INIT[2164], INIT[1652], INIT[1140], INIT[ 628], INIT[ 116],
  INIT[3699], INIT[3187], INIT[2675], INIT[2163], INIT[1651], INIT[1139], INIT[ 627], INIT[ 115],
  INIT[3698], INIT[3186], INIT[2674], INIT[2162], INIT[1650], INIT[1138], INIT[ 626], INIT[ 114],
  INIT[3697], INIT[3185], INIT[2673], INIT[2161], INIT[1649], INIT[1137], INIT[ 625], INIT[ 113],
  INIT[3696], INIT[3184], INIT[2672], INIT[2160], INIT[1648], INIT[1136], INIT[ 624], INIT[ 112],
  INIT[3695], INIT[3183], INIT[2671], INIT[2159], INIT[1647], INIT[1135], INIT[ 623], INIT[ 111],
  INIT[3694], INIT[3182], INIT[2670], INIT[2158], INIT[1646], INIT[1134], INIT[ 622], INIT[ 110],
  INIT[3693], INIT[3181], INIT[2669], INIT[2157], INIT[1645], INIT[1133], INIT[ 621], INIT[ 109],
  INIT[3692], INIT[3180], INIT[2668], INIT[2156], INIT[1644], INIT[1132], INIT[ 620], INIT[ 108],
  INIT[3691], INIT[3179], INIT[2667], INIT[2155], INIT[1643], INIT[1131], INIT[ 619], INIT[ 107],
  INIT[3690], INIT[3178], INIT[2666], INIT[2154], INIT[1642], INIT[1130], INIT[ 618], INIT[ 106],
  INIT[3689], INIT[3177], INIT[2665], INIT[2153], INIT[1641], INIT[1129], INIT[ 617], INIT[ 105],
  INIT[3688], INIT[3176], INIT[2664], INIT[2152], INIT[1640], INIT[1128], INIT[ 616], INIT[ 104],
  INIT[3687], INIT[3175], INIT[2663], INIT[2151], INIT[1639], INIT[1127], INIT[ 615], INIT[ 103],
  INIT[3686], INIT[3174], INIT[2662], INIT[2150], INIT[1638], INIT[1126], INIT[ 614], INIT[ 102],
  INIT[3685], INIT[3173], INIT[2661], INIT[2149], INIT[1637], INIT[1125], INIT[ 613], INIT[ 101],
  INIT[3684], INIT[3172], INIT[2660], INIT[2148], INIT[1636], INIT[1124], INIT[ 612], INIT[ 100],
  INIT[3683], INIT[3171], INIT[2659], INIT[2147], INIT[1635], INIT[1123], INIT[ 611], INIT[  99],
  INIT[3682], INIT[3170], INIT[2658], INIT[2146], INIT[1634], INIT[1122], INIT[ 610], INIT[  98],
  INIT[3681], INIT[3169], INIT[2657], INIT[2145], INIT[1633], INIT[1121], INIT[ 609], INIT[  97],
  INIT[3680], INIT[3168], INIT[2656], INIT[2144], INIT[1632], INIT[1120], INIT[ 608], INIT[  96]
};
localparam [255:0] INIT_4 = {
  INIT[3743], INIT[3231], INIT[2719], INIT[2207], INIT[1695], INIT[1183], INIT[ 671], INIT[ 159],
  INIT[3742], INIT[3230], INIT[2718], INIT[2206], INIT[1694], INIT[1182], INIT[ 670], INIT[ 158],
  INIT[3741], INIT[3229], INIT[2717], INIT[2205], INIT[1693], INIT[1181], INIT[ 669], INIT[ 157],
  INIT[3740], INIT[3228], INIT[2716], INIT[2204], INIT[1692], INIT[1180], INIT[ 668], INIT[ 156],
  INIT[3739], INIT[3227], INIT[2715], INIT[2203], INIT[1691], INIT[1179], INIT[ 667], INIT[ 155],
  INIT[3738], INIT[3226], INIT[2714], INIT[2202], INIT[1690], INIT[1178], INIT[ 666], INIT[ 154],
  INIT[3737], INIT[3225], INIT[2713], INIT[2201], INIT[1689], INIT[1177], INIT[ 665], INIT[ 153],
  INIT[3736], INIT[3224], INIT[2712], INIT[2200], INIT[1688], INIT[1176], INIT[ 664], INIT[ 152],
  INIT[3735], INIT[3223], INIT[2711], INIT[2199], INIT[1687], INIT[1175], INIT[ 663], INIT[ 151],
  INIT[3734], INIT[3222], INIT[2710], INIT[2198], INIT[1686], INIT[1174], INIT[ 662], INIT[ 150],
  INIT[3733], INIT[3221], INIT[2709], INIT[2197], INIT[1685], INIT[1173], INIT[ 661], INIT[ 149],
  INIT[3732], INIT[3220], INIT[2708], INIT[2196], INIT[1684], INIT[1172], INIT[ 660], INIT[ 148],
  INIT[3731], INIT[3219], INIT[2707], INIT[2195], INIT[1683], INIT[1171], INIT[ 659], INIT[ 147],
  INIT[3730], INIT[3218], INIT[2706], INIT[2194], INIT[1682], INIT[1170], INIT[ 658], INIT[ 146],
  INIT[3729], INIT[3217], INIT[2705], INIT[2193], INIT[1681], INIT[1169], INIT[ 657], INIT[ 145],
  INIT[3728], INIT[3216], INIT[2704], INIT[2192], INIT[1680], INIT[1168], INIT[ 656], INIT[ 144],
  INIT[3727], INIT[3215], INIT[2703], INIT[2191], INIT[1679], INIT[1167], INIT[ 655], INIT[ 143],
  INIT[3726], INIT[3214], INIT[2702], INIT[2190], INIT[1678], INIT[1166], INIT[ 654], INIT[ 142],
  INIT[3725], INIT[3213], INIT[2701], INIT[2189], INIT[1677], INIT[1165], INIT[ 653], INIT[ 141],
  INIT[3724], INIT[3212], INIT[2700], INIT[2188], INIT[1676], INIT[1164], INIT[ 652], INIT[ 140],
  INIT[3723], INIT[3211], INIT[2699], INIT[2187], INIT[1675], INIT[1163], INIT[ 651], INIT[ 139],
  INIT[3722], INIT[3210], INIT[2698], INIT[2186], INIT[1674], INIT[1162], INIT[ 650], INIT[ 138],
  INIT[3721], INIT[3209], INIT[2697], INIT[2185], INIT[1673], INIT[1161], INIT[ 649], INIT[ 137],
  INIT[3720], INIT[3208], INIT[2696], INIT[2184], INIT[1672], INIT[1160], INIT[ 648], INIT[ 136],
  INIT[3719], INIT[3207], INIT[2695], INIT[2183], INIT[1671], INIT[1159], INIT[ 647], INIT[ 135],
  INIT[3718], INIT[3206], INIT[2694], INIT[2182], INIT[1670], INIT[1158], INIT[ 646], INIT[ 134],
  INIT[3717], INIT[3205], INIT[2693], INIT[2181], INIT[1669], INIT[1157], INIT[ 645], INIT[ 133],
  INIT[3716], INIT[3204], INIT[2692], INIT[2180], INIT[1668], INIT[1156], INIT[ 644], INIT[ 132],
  INIT[3715], INIT[3203], INIT[2691], INIT[2179], INIT[1667], INIT[1155], INIT[ 643], INIT[ 131],
  INIT[3714], INIT[3202], INIT[2690], INIT[2178], INIT[1666], INIT[1154], INIT[ 642], INIT[ 130],
  INIT[3713], INIT[3201], INIT[2689], INIT[2177], INIT[1665], INIT[1153], INIT[ 641], INIT[ 129],
  INIT[3712], INIT[3200], INIT[2688], INIT[2176], INIT[1664], INIT[1152], INIT[ 640], INIT[ 128]
};
localparam [255:0] INIT_5 = {
  INIT[3775], INIT[3263], INIT[2751], INIT[2239], INIT[1727], INIT[1215], INIT[ 703], INIT[ 191],
  INIT[3774], INIT[3262], INIT[2750], INIT[2238], INIT[1726], INIT[1214], INIT[ 702], INIT[ 190],
  INIT[3773], INIT[3261], INIT[2749], INIT[2237], INIT[1725], INIT[1213], INIT[ 701], INIT[ 189],
  INIT[3772], INIT[3260], INIT[2748], INIT[2236], INIT[1724], INIT[1212], INIT[ 700], INIT[ 188],
  INIT[3771], INIT[3259], INIT[2747], INIT[2235], INIT[1723], INIT[1211], INIT[ 699], INIT[ 187],
  INIT[3770], INIT[3258], INIT[2746], INIT[2234], INIT[1722], INIT[1210], INIT[ 698], INIT[ 186],
  INIT[3769], INIT[3257], INIT[2745], INIT[2233], INIT[1721], INIT[1209], INIT[ 697], INIT[ 185],
  INIT[3768], INIT[3256], INIT[2744], INIT[2232], INIT[1720], INIT[1208], INIT[ 696], INIT[ 184],
  INIT[3767], INIT[3255], INIT[2743], INIT[2231], INIT[1719], INIT[1207], INIT[ 695], INIT[ 183],
  INIT[3766], INIT[3254], INIT[2742], INIT[2230], INIT[1718], INIT[1206], INIT[ 694], INIT[ 182],
  INIT[3765], INIT[3253], INIT[2741], INIT[2229], INIT[1717], INIT[1205], INIT[ 693], INIT[ 181],
  INIT[3764], INIT[3252], INIT[2740], INIT[2228], INIT[1716], INIT[1204], INIT[ 692], INIT[ 180],
  INIT[3763], INIT[3251], INIT[2739], INIT[2227], INIT[1715], INIT[1203], INIT[ 691], INIT[ 179],
  INIT[3762], INIT[3250], INIT[2738], INIT[2226], INIT[1714], INIT[1202], INIT[ 690], INIT[ 178],
  INIT[3761], INIT[3249], INIT[2737], INIT[2225], INIT[1713], INIT[1201], INIT[ 689], INIT[ 177],
  INIT[3760], INIT[3248], INIT[2736], INIT[2224], INIT[1712], INIT[1200], INIT[ 688], INIT[ 176],
  INIT[3759], INIT[3247], INIT[2735], INIT[2223], INIT[1711], INIT[1199], INIT[ 687], INIT[ 175],
  INIT[3758], INIT[3246], INIT[2734], INIT[2222], INIT[1710], INIT[1198], INIT[ 686], INIT[ 174],
  INIT[3757], INIT[3245], INIT[2733], INIT[2221], INIT[1709], INIT[1197], INIT[ 685], INIT[ 173],
  INIT[3756], INIT[3244], INIT[2732], INIT[2220], INIT[1708], INIT[1196], INIT[ 684], INIT[ 172],
  INIT[3755], INIT[3243], INIT[2731], INIT[2219], INIT[1707], INIT[1195], INIT[ 683], INIT[ 171],
  INIT[3754], INIT[3242], INIT[2730], INIT[2218], INIT[1706], INIT[1194], INIT[ 682], INIT[ 170],
  INIT[3753], INIT[3241], INIT[2729], INIT[2217], INIT[1705], INIT[1193], INIT[ 681], INIT[ 169],
  INIT[3752], INIT[3240], INIT[2728], INIT[2216], INIT[1704], INIT[1192], INIT[ 680], INIT[ 168],
  INIT[3751], INIT[3239], INIT[2727], INIT[2215], INIT[1703], INIT[1191], INIT[ 679], INIT[ 167],
  INIT[3750], INIT[3238], INIT[2726], INIT[2214], INIT[1702], INIT[1190], INIT[ 678], INIT[ 166],
  INIT[3749], INIT[3237], INIT[2725], INIT[2213], INIT[1701], INIT[1189], INIT[ 677], INIT[ 165],
  INIT[3748], INIT[3236], INIT[2724], INIT[2212], INIT[1700], INIT[1188], INIT[ 676], INIT[ 164],
  INIT[3747], INIT[3235], INIT[2723], INIT[2211], INIT[1699], INIT[1187], INIT[ 675], INIT[ 163],
  INIT[3746], INIT[3234], INIT[2722], INIT[2210], INIT[1698], INIT[1186], INIT[ 674], INIT[ 162],
  INIT[3745], INIT[3233], INIT[2721], INIT[2209], INIT[1697], INIT[1185], INIT[ 673], INIT[ 161],
  INIT[3744], INIT[3232], INIT[2720], INIT[2208], INIT[1696], INIT[1184], INIT[ 672], INIT[ 160]
};
localparam [255:0] INIT_6 = {
  INIT[3807], INIT[3295], INIT[2783], INIT[2271], INIT[1759], INIT[1247], INIT[ 735], INIT[ 223],
  INIT[3806], INIT[3294], INIT[2782], INIT[2270], INIT[1758], INIT[1246], INIT[ 734], INIT[ 222],
  INIT[3805], INIT[3293], INIT[2781], INIT[2269], INIT[1757], INIT[1245], INIT[ 733], INIT[ 221],
  INIT[3804], INIT[3292], INIT[2780], INIT[2268], INIT[1756], INIT[1244], INIT[ 732], INIT[ 220],
  INIT[3803], INIT[3291], INIT[2779], INIT[2267], INIT[1755], INIT[1243], INIT[ 731], INIT[ 219],
  INIT[3802], INIT[3290], INIT[2778], INIT[2266], INIT[1754], INIT[1242], INIT[ 730], INIT[ 218],
  INIT[3801], INIT[3289], INIT[2777], INIT[2265], INIT[1753], INIT[1241], INIT[ 729], INIT[ 217],
  INIT[3800], INIT[3288], INIT[2776], INIT[2264], INIT[1752], INIT[1240], INIT[ 728], INIT[ 216],
  INIT[3799], INIT[3287], INIT[2775], INIT[2263], INIT[1751], INIT[1239], INIT[ 727], INIT[ 215],
  INIT[3798], INIT[3286], INIT[2774], INIT[2262], INIT[1750], INIT[1238], INIT[ 726], INIT[ 214],
  INIT[3797], INIT[3285], INIT[2773], INIT[2261], INIT[1749], INIT[1237], INIT[ 725], INIT[ 213],
  INIT[3796], INIT[3284], INIT[2772], INIT[2260], INIT[1748], INIT[1236], INIT[ 724], INIT[ 212],
  INIT[3795], INIT[3283], INIT[2771], INIT[2259], INIT[1747], INIT[1235], INIT[ 723], INIT[ 211],
  INIT[3794], INIT[3282], INIT[2770], INIT[2258], INIT[1746], INIT[1234], INIT[ 722], INIT[ 210],
  INIT[3793], INIT[3281], INIT[2769], INIT[2257], INIT[1745], INIT[1233], INIT[ 721], INIT[ 209],
  INIT[3792], INIT[3280], INIT[2768], INIT[2256], INIT[1744], INIT[1232], INIT[ 720], INIT[ 208],
  INIT[3791], INIT[3279], INIT[2767], INIT[2255], INIT[1743], INIT[1231], INIT[ 719], INIT[ 207],
  INIT[3790], INIT[3278], INIT[2766], INIT[2254], INIT[1742], INIT[1230], INIT[ 718], INIT[ 206],
  INIT[3789], INIT[3277], INIT[2765], INIT[2253], INIT[1741], INIT[1229], INIT[ 717], INIT[ 205],
  INIT[3788], INIT[3276], INIT[2764], INIT[2252], INIT[1740], INIT[1228], INIT[ 716], INIT[ 204],
  INIT[3787], INIT[3275], INIT[2763], INIT[2251], INIT[1739], INIT[1227], INIT[ 715], INIT[ 203],
  INIT[3786], INIT[3274], INIT[2762], INIT[2250], INIT[1738], INIT[1226], INIT[ 714], INIT[ 202],
  INIT[3785], INIT[3273], INIT[2761], INIT[2249], INIT[1737], INIT[1225], INIT[ 713], INIT[ 201],
  INIT[3784], INIT[3272], INIT[2760], INIT[2248], INIT[1736], INIT[1224], INIT[ 712], INIT[ 200],
  INIT[3783], INIT[3271], INIT[2759], INIT[2247], INIT[1735], INIT[1223], INIT[ 711], INIT[ 199],
  INIT[3782], INIT[3270], INIT[2758], INIT[2246], INIT[1734], INIT[1222], INIT[ 710], INIT[ 198],
  INIT[3781], INIT[3269], INIT[2757], INIT[2245], INIT[1733], INIT[1221], INIT[ 709], INIT[ 197],
  INIT[3780], INIT[3268], INIT[2756], INIT[2244], INIT[1732], INIT[1220], INIT[ 708], INIT[ 196],
  INIT[3779], INIT[3267], INIT[2755], INIT[2243], INIT[1731], INIT[1219], INIT[ 707], INIT[ 195],
  INIT[3778], INIT[3266], INIT[2754], INIT[2242], INIT[1730], INIT[1218], INIT[ 706], INIT[ 194],
  INIT[3777], INIT[3265], INIT[2753], INIT[2241], INIT[1729], INIT[1217], INIT[ 705], INIT[ 193],
  INIT[3776], INIT[3264], INIT[2752], INIT[2240], INIT[1728], INIT[1216], INIT[ 704], INIT[ 192]
};
localparam [255:0] INIT_7 = {
  INIT[3839], INIT[3327], INIT[2815], INIT[2303], INIT[1791], INIT[1279], INIT[ 767], INIT[ 255],
  INIT[3838], INIT[3326], INIT[2814], INIT[2302], INIT[1790], INIT[1278], INIT[ 766], INIT[ 254],
  INIT[3837], INIT[3325], INIT[2813], INIT[2301], INIT[1789], INIT[1277], INIT[ 765], INIT[ 253],
  INIT[3836], INIT[3324], INIT[2812], INIT[2300], INIT[1788], INIT[1276], INIT[ 764], INIT[ 252],
  INIT[3835], INIT[3323], INIT[2811], INIT[2299], INIT[1787], INIT[1275], INIT[ 763], INIT[ 251],
  INIT[3834], INIT[3322], INIT[2810], INIT[2298], INIT[1786], INIT[1274], INIT[ 762], INIT[ 250],
  INIT[3833], INIT[3321], INIT[2809], INIT[2297], INIT[1785], INIT[1273], INIT[ 761], INIT[ 249],
  INIT[3832], INIT[3320], INIT[2808], INIT[2296], INIT[1784], INIT[1272], INIT[ 760], INIT[ 248],
  INIT[3831], INIT[3319], INIT[2807], INIT[2295], INIT[1783], INIT[1271], INIT[ 759], INIT[ 247],
  INIT[3830], INIT[3318], INIT[2806], INIT[2294], INIT[1782], INIT[1270], INIT[ 758], INIT[ 246],
  INIT[3829], INIT[3317], INIT[2805], INIT[2293], INIT[1781], INIT[1269], INIT[ 757], INIT[ 245],
  INIT[3828], INIT[3316], INIT[2804], INIT[2292], INIT[1780], INIT[1268], INIT[ 756], INIT[ 244],
  INIT[3827], INIT[3315], INIT[2803], INIT[2291], INIT[1779], INIT[1267], INIT[ 755], INIT[ 243],
  INIT[3826], INIT[3314], INIT[2802], INIT[2290], INIT[1778], INIT[1266], INIT[ 754], INIT[ 242],
  INIT[3825], INIT[3313], INIT[2801], INIT[2289], INIT[1777], INIT[1265], INIT[ 753], INIT[ 241],
  INIT[3824], INIT[3312], INIT[2800], INIT[2288], INIT[1776], INIT[1264], INIT[ 752], INIT[ 240],
  INIT[3823], INIT[3311], INIT[2799], INIT[2287], INIT[1775], INIT[1263], INIT[ 751], INIT[ 239],
  INIT[3822], INIT[3310], INIT[2798], INIT[2286], INIT[1774], INIT[1262], INIT[ 750], INIT[ 238],
  INIT[3821], INIT[3309], INIT[2797], INIT[2285], INIT[1773], INIT[1261], INIT[ 749], INIT[ 237],
  INIT[3820], INIT[3308], INIT[2796], INIT[2284], INIT[1772], INIT[1260], INIT[ 748], INIT[ 236],
  INIT[3819], INIT[3307], INIT[2795], INIT[2283], INIT[1771], INIT[1259], INIT[ 747], INIT[ 235],
  INIT[3818], INIT[3306], INIT[2794], INIT[2282], INIT[1770], INIT[1258], INIT[ 746], INIT[ 234],
  INIT[3817], INIT[3305], INIT[2793], INIT[2281], INIT[1769], INIT[1257], INIT[ 745], INIT[ 233],
  INIT[3816], INIT[3304], INIT[2792], INIT[2280], INIT[1768], INIT[1256], INIT[ 744], INIT[ 232],
  INIT[3815], INIT[3303], INIT[2791], INIT[2279], INIT[1767], INIT[1255], INIT[ 743], INIT[ 231],
  INIT[3814], INIT[3302], INIT[2790], INIT[2278], INIT[1766], INIT[1254], INIT[ 742], INIT[ 230],
  INIT[3813], INIT[3301], INIT[2789], INIT[2277], INIT[1765], INIT[1253], INIT[ 741], INIT[ 229],
  INIT[3812], INIT[3300], INIT[2788], INIT[2276], INIT[1764], INIT[1252], INIT[ 740], INIT[ 228],
  INIT[3811], INIT[3299], INIT[2787], INIT[2275], INIT[1763], INIT[1251], INIT[ 739], INIT[ 227],
  INIT[3810], INIT[3298], INIT[2786], INIT[2274], INIT[1762], INIT[1250], INIT[ 738], INIT[ 226],
  INIT[3809], INIT[3297], INIT[2785], INIT[2273], INIT[1761], INIT[1249], INIT[ 737], INIT[ 225],
  INIT[3808], INIT[3296], INIT[2784], INIT[2272], INIT[1760], INIT[1248], INIT[ 736], INIT[ 224]
};
localparam [255:0] INIT_8 = {
  INIT[3871], INIT[3359], INIT[2847], INIT[2335], INIT[1823], INIT[1311], INIT[ 799], INIT[ 287],
  INIT[3870], INIT[3358], INIT[2846], INIT[2334], INIT[1822], INIT[1310], INIT[ 798], INIT[ 286],
  INIT[3869], INIT[3357], INIT[2845], INIT[2333], INIT[1821], INIT[1309], INIT[ 797], INIT[ 285],
  INIT[3868], INIT[3356], INIT[2844], INIT[2332], INIT[1820], INIT[1308], INIT[ 796], INIT[ 284],
  INIT[3867], INIT[3355], INIT[2843], INIT[2331], INIT[1819], INIT[1307], INIT[ 795], INIT[ 283],
  INIT[3866], INIT[3354], INIT[2842], INIT[2330], INIT[1818], INIT[1306], INIT[ 794], INIT[ 282],
  INIT[3865], INIT[3353], INIT[2841], INIT[2329], INIT[1817], INIT[1305], INIT[ 793], INIT[ 281],
  INIT[3864], INIT[3352], INIT[2840], INIT[2328], INIT[1816], INIT[1304], INIT[ 792], INIT[ 280],
  INIT[3863], INIT[3351], INIT[2839], INIT[2327], INIT[1815], INIT[1303], INIT[ 791], INIT[ 279],
  INIT[3862], INIT[3350], INIT[2838], INIT[2326], INIT[1814], INIT[1302], INIT[ 790], INIT[ 278],
  INIT[3861], INIT[3349], INIT[2837], INIT[2325], INIT[1813], INIT[1301], INIT[ 789], INIT[ 277],
  INIT[3860], INIT[3348], INIT[2836], INIT[2324], INIT[1812], INIT[1300], INIT[ 788], INIT[ 276],
  INIT[3859], INIT[3347], INIT[2835], INIT[2323], INIT[1811], INIT[1299], INIT[ 787], INIT[ 275],
  INIT[3858], INIT[3346], INIT[2834], INIT[2322], INIT[1810], INIT[1298], INIT[ 786], INIT[ 274],
  INIT[3857], INIT[3345], INIT[2833], INIT[2321], INIT[1809], INIT[1297], INIT[ 785], INIT[ 273],
  INIT[3856], INIT[3344], INIT[2832], INIT[2320], INIT[1808], INIT[1296], INIT[ 784], INIT[ 272],
  INIT[3855], INIT[3343], INIT[2831], INIT[2319], INIT[1807], INIT[1295], INIT[ 783], INIT[ 271],
  INIT[3854], INIT[3342], INIT[2830], INIT[2318], INIT[1806], INIT[1294], INIT[ 782], INIT[ 270],
  INIT[3853], INIT[3341], INIT[2829], INIT[2317], INIT[1805], INIT[1293], INIT[ 781], INIT[ 269],
  INIT[3852], INIT[3340], INIT[2828], INIT[2316], INIT[1804], INIT[1292], INIT[ 780], INIT[ 268],
  INIT[3851], INIT[3339], INIT[2827], INIT[2315], INIT[1803], INIT[1291], INIT[ 779], INIT[ 267],
  INIT[3850], INIT[3338], INIT[2826], INIT[2314], INIT[1802], INIT[1290], INIT[ 778], INIT[ 266],
  INIT[3849], INIT[3337], INIT[2825], INIT[2313], INIT[1801], INIT[1289], INIT[ 777], INIT[ 265],
  INIT[3848], INIT[3336], INIT[2824], INIT[2312], INIT[1800], INIT[1288], INIT[ 776], INIT[ 264],
  INIT[3847], INIT[3335], INIT[2823], INIT[2311], INIT[1799], INIT[1287], INIT[ 775], INIT[ 263],
  INIT[3846], INIT[3334], INIT[2822], INIT[2310], INIT[1798], INIT[1286], INIT[ 774], INIT[ 262],
  INIT[3845], INIT[3333], INIT[2821], INIT[2309], INIT[1797], INIT[1285], INIT[ 773], INIT[ 261],
  INIT[3844], INIT[3332], INIT[2820], INIT[2308], INIT[1796], INIT[1284], INIT[ 772], INIT[ 260],
  INIT[3843], INIT[3331], INIT[2819], INIT[2307], INIT[1795], INIT[1283], INIT[ 771], INIT[ 259],
  INIT[3842], INIT[3330], INIT[2818], INIT[2306], INIT[1794], INIT[1282], INIT[ 770], INIT[ 258],
  INIT[3841], INIT[3329], INIT[2817], INIT[2305], INIT[1793], INIT[1281], INIT[ 769], INIT[ 257],
  INIT[3840], INIT[3328], INIT[2816], INIT[2304], INIT[1792], INIT[1280], INIT[ 768], INIT[ 256]
};
localparam [255:0] INIT_9 = {
  INIT[3903], INIT[3391], INIT[2879], INIT[2367], INIT[1855], INIT[1343], INIT[ 831], INIT[ 319],
  INIT[3902], INIT[3390], INIT[2878], INIT[2366], INIT[1854], INIT[1342], INIT[ 830], INIT[ 318],
  INIT[3901], INIT[3389], INIT[2877], INIT[2365], INIT[1853], INIT[1341], INIT[ 829], INIT[ 317],
  INIT[3900], INIT[3388], INIT[2876], INIT[2364], INIT[1852], INIT[1340], INIT[ 828], INIT[ 316],
  INIT[3899], INIT[3387], INIT[2875], INIT[2363], INIT[1851], INIT[1339], INIT[ 827], INIT[ 315],
  INIT[3898], INIT[3386], INIT[2874], INIT[2362], INIT[1850], INIT[1338], INIT[ 826], INIT[ 314],
  INIT[3897], INIT[3385], INIT[2873], INIT[2361], INIT[1849], INIT[1337], INIT[ 825], INIT[ 313],
  INIT[3896], INIT[3384], INIT[2872], INIT[2360], INIT[1848], INIT[1336], INIT[ 824], INIT[ 312],
  INIT[3895], INIT[3383], INIT[2871], INIT[2359], INIT[1847], INIT[1335], INIT[ 823], INIT[ 311],
  INIT[3894], INIT[3382], INIT[2870], INIT[2358], INIT[1846], INIT[1334], INIT[ 822], INIT[ 310],
  INIT[3893], INIT[3381], INIT[2869], INIT[2357], INIT[1845], INIT[1333], INIT[ 821], INIT[ 309],
  INIT[3892], INIT[3380], INIT[2868], INIT[2356], INIT[1844], INIT[1332], INIT[ 820], INIT[ 308],
  INIT[3891], INIT[3379], INIT[2867], INIT[2355], INIT[1843], INIT[1331], INIT[ 819], INIT[ 307],
  INIT[3890], INIT[3378], INIT[2866], INIT[2354], INIT[1842], INIT[1330], INIT[ 818], INIT[ 306],
  INIT[3889], INIT[3377], INIT[2865], INIT[2353], INIT[1841], INIT[1329], INIT[ 817], INIT[ 305],
  INIT[3888], INIT[3376], INIT[2864], INIT[2352], INIT[1840], INIT[1328], INIT[ 816], INIT[ 304],
  INIT[3887], INIT[3375], INIT[2863], INIT[2351], INIT[1839], INIT[1327], INIT[ 815], INIT[ 303],
  INIT[3886], INIT[3374], INIT[2862], INIT[2350], INIT[1838], INIT[1326], INIT[ 814], INIT[ 302],
  INIT[3885], INIT[3373], INIT[2861], INIT[2349], INIT[1837], INIT[1325], INIT[ 813], INIT[ 301],
  INIT[3884], INIT[3372], INIT[2860], INIT[2348], INIT[1836], INIT[1324], INIT[ 812], INIT[ 300],
  INIT[3883], INIT[3371], INIT[2859], INIT[2347], INIT[1835], INIT[1323], INIT[ 811], INIT[ 299],
  INIT[3882], INIT[3370], INIT[2858], INIT[2346], INIT[1834], INIT[1322], INIT[ 810], INIT[ 298],
  INIT[3881], INIT[3369], INIT[2857], INIT[2345], INIT[1833], INIT[1321], INIT[ 809], INIT[ 297],
  INIT[3880], INIT[3368], INIT[2856], INIT[2344], INIT[1832], INIT[1320], INIT[ 808], INIT[ 296],
  INIT[3879], INIT[3367], INIT[2855], INIT[2343], INIT[1831], INIT[1319], INIT[ 807], INIT[ 295],
  INIT[3878], INIT[3366], INIT[2854], INIT[2342], INIT[1830], INIT[1318], INIT[ 806], INIT[ 294],
  INIT[3877], INIT[3365], INIT[2853], INIT[2341], INIT[1829], INIT[1317], INIT[ 805], INIT[ 293],
  INIT[3876], INIT[3364], INIT[2852], INIT[2340], INIT[1828], INIT[1316], INIT[ 804], INIT[ 292],
  INIT[3875], INIT[3363], INIT[2851], INIT[2339], INIT[1827], INIT[1315], INIT[ 803], INIT[ 291],
  INIT[3874], INIT[3362], INIT[2850], INIT[2338], INIT[1826], INIT[1314], INIT[ 802], INIT[ 290],
  INIT[3873], INIT[3361], INIT[2849], INIT[2337], INIT[1825], INIT[1313], INIT[ 801], INIT[ 289],
  INIT[3872], INIT[3360], INIT[2848], INIT[2336], INIT[1824], INIT[1312], INIT[ 800], INIT[ 288]
};
localparam [255:0] INIT_A = {
  INIT[3935], INIT[3423], INIT[2911], INIT[2399], INIT[1887], INIT[1375], INIT[ 863], INIT[ 351],
  INIT[3934], INIT[3422], INIT[2910], INIT[2398], INIT[1886], INIT[1374], INIT[ 862], INIT[ 350],
  INIT[3933], INIT[3421], INIT[2909], INIT[2397], INIT[1885], INIT[1373], INIT[ 861], INIT[ 349],
  INIT[3932], INIT[3420], INIT[2908], INIT[2396], INIT[1884], INIT[1372], INIT[ 860], INIT[ 348],
  INIT[3931], INIT[3419], INIT[2907], INIT[2395], INIT[1883], INIT[1371], INIT[ 859], INIT[ 347],
  INIT[3930], INIT[3418], INIT[2906], INIT[2394], INIT[1882], INIT[1370], INIT[ 858], INIT[ 346],
  INIT[3929], INIT[3417], INIT[2905], INIT[2393], INIT[1881], INIT[1369], INIT[ 857], INIT[ 345],
  INIT[3928], INIT[3416], INIT[2904], INIT[2392], INIT[1880], INIT[1368], INIT[ 856], INIT[ 344],
  INIT[3927], INIT[3415], INIT[2903], INIT[2391], INIT[1879], INIT[1367], INIT[ 855], INIT[ 343],
  INIT[3926], INIT[3414], INIT[2902], INIT[2390], INIT[1878], INIT[1366], INIT[ 854], INIT[ 342],
  INIT[3925], INIT[3413], INIT[2901], INIT[2389], INIT[1877], INIT[1365], INIT[ 853], INIT[ 341],
  INIT[3924], INIT[3412], INIT[2900], INIT[2388], INIT[1876], INIT[1364], INIT[ 852], INIT[ 340],
  INIT[3923], INIT[3411], INIT[2899], INIT[2387], INIT[1875], INIT[1363], INIT[ 851], INIT[ 339],
  INIT[3922], INIT[3410], INIT[2898], INIT[2386], INIT[1874], INIT[1362], INIT[ 850], INIT[ 338],
  INIT[3921], INIT[3409], INIT[2897], INIT[2385], INIT[1873], INIT[1361], INIT[ 849], INIT[ 337],
  INIT[3920], INIT[3408], INIT[2896], INIT[2384], INIT[1872], INIT[1360], INIT[ 848], INIT[ 336],
  INIT[3919], INIT[3407], INIT[2895], INIT[2383], INIT[1871], INIT[1359], INIT[ 847], INIT[ 335],
  INIT[3918], INIT[3406], INIT[2894], INIT[2382], INIT[1870], INIT[1358], INIT[ 846], INIT[ 334],
  INIT[3917], INIT[3405], INIT[2893], INIT[2381], INIT[1869], INIT[1357], INIT[ 845], INIT[ 333],
  INIT[3916], INIT[3404], INIT[2892], INIT[2380], INIT[1868], INIT[1356], INIT[ 844], INIT[ 332],
  INIT[3915], INIT[3403], INIT[2891], INIT[2379], INIT[1867], INIT[1355], INIT[ 843], INIT[ 331],
  INIT[3914], INIT[3402], INIT[2890], INIT[2378], INIT[1866], INIT[1354], INIT[ 842], INIT[ 330],
  INIT[3913], INIT[3401], INIT[2889], INIT[2377], INIT[1865], INIT[1353], INIT[ 841], INIT[ 329],
  INIT[3912], INIT[3400], INIT[2888], INIT[2376], INIT[1864], INIT[1352], INIT[ 840], INIT[ 328],
  INIT[3911], INIT[3399], INIT[2887], INIT[2375], INIT[1863], INIT[1351], INIT[ 839], INIT[ 327],
  INIT[3910], INIT[3398], INIT[2886], INIT[2374], INIT[1862], INIT[1350], INIT[ 838], INIT[ 326],
  INIT[3909], INIT[3397], INIT[2885], INIT[2373], INIT[1861], INIT[1349], INIT[ 837], INIT[ 325],
  INIT[3908], INIT[3396], INIT[2884], INIT[2372], INIT[1860], INIT[1348], INIT[ 836], INIT[ 324],
  INIT[3907], INIT[3395], INIT[2883], INIT[2371], INIT[1859], INIT[1347], INIT[ 835], INIT[ 323],
  INIT[3906], INIT[3394], INIT[2882], INIT[2370], INIT[1858], INIT[1346], INIT[ 834], INIT[ 322],
  INIT[3905], INIT[3393], INIT[2881], INIT[2369], INIT[1857], INIT[1345], INIT[ 833], INIT[ 321],
  INIT[3904], INIT[3392], INIT[2880], INIT[2368], INIT[1856], INIT[1344], INIT[ 832], INIT[ 320]
};
localparam [255:0] INIT_B = {
  INIT[3967], INIT[3455], INIT[2943], INIT[2431], INIT[1919], INIT[1407], INIT[ 895], INIT[ 383],
  INIT[3966], INIT[3454], INIT[2942], INIT[2430], INIT[1918], INIT[1406], INIT[ 894], INIT[ 382],
  INIT[3965], INIT[3453], INIT[2941], INIT[2429], INIT[1917], INIT[1405], INIT[ 893], INIT[ 381],
  INIT[3964], INIT[3452], INIT[2940], INIT[2428], INIT[1916], INIT[1404], INIT[ 892], INIT[ 380],
  INIT[3963], INIT[3451], INIT[2939], INIT[2427], INIT[1915], INIT[1403], INIT[ 891], INIT[ 379],
  INIT[3962], INIT[3450], INIT[2938], INIT[2426], INIT[1914], INIT[1402], INIT[ 890], INIT[ 378],
  INIT[3961], INIT[3449], INIT[2937], INIT[2425], INIT[1913], INIT[1401], INIT[ 889], INIT[ 377],
  INIT[3960], INIT[3448], INIT[2936], INIT[2424], INIT[1912], INIT[1400], INIT[ 888], INIT[ 376],
  INIT[3959], INIT[3447], INIT[2935], INIT[2423], INIT[1911], INIT[1399], INIT[ 887], INIT[ 375],
  INIT[3958], INIT[3446], INIT[2934], INIT[2422], INIT[1910], INIT[1398], INIT[ 886], INIT[ 374],
  INIT[3957], INIT[3445], INIT[2933], INIT[2421], INIT[1909], INIT[1397], INIT[ 885], INIT[ 373],
  INIT[3956], INIT[3444], INIT[2932], INIT[2420], INIT[1908], INIT[1396], INIT[ 884], INIT[ 372],
  INIT[3955], INIT[3443], INIT[2931], INIT[2419], INIT[1907], INIT[1395], INIT[ 883], INIT[ 371],
  INIT[3954], INIT[3442], INIT[2930], INIT[2418], INIT[1906], INIT[1394], INIT[ 882], INIT[ 370],
  INIT[3953], INIT[3441], INIT[2929], INIT[2417], INIT[1905], INIT[1393], INIT[ 881], INIT[ 369],
  INIT[3952], INIT[3440], INIT[2928], INIT[2416], INIT[1904], INIT[1392], INIT[ 880], INIT[ 368],
  INIT[3951], INIT[3439], INIT[2927], INIT[2415], INIT[1903], INIT[1391], INIT[ 879], INIT[ 367],
  INIT[3950], INIT[3438], INIT[2926], INIT[2414], INIT[1902], INIT[1390], INIT[ 878], INIT[ 366],
  INIT[3949], INIT[3437], INIT[2925], INIT[2413], INIT[1901], INIT[1389], INIT[ 877], INIT[ 365],
  INIT[3948], INIT[3436], INIT[2924], INIT[2412], INIT[1900], INIT[1388], INIT[ 876], INIT[ 364],
  INIT[3947], INIT[3435], INIT[2923], INIT[2411], INIT[1899], INIT[1387], INIT[ 875], INIT[ 363],
  INIT[3946], INIT[3434], INIT[2922], INIT[2410], INIT[1898], INIT[1386], INIT[ 874], INIT[ 362],
  INIT[3945], INIT[3433], INIT[2921], INIT[2409], INIT[1897], INIT[1385], INIT[ 873], INIT[ 361],
  INIT[3944], INIT[3432], INIT[2920], INIT[2408], INIT[1896], INIT[1384], INIT[ 872], INIT[ 360],
  INIT[3943], INIT[3431], INIT[2919], INIT[2407], INIT[1895], INIT[1383], INIT[ 871], INIT[ 359],
  INIT[3942], INIT[3430], INIT[2918], INIT[2406], INIT[1894], INIT[1382], INIT[ 870], INIT[ 358],
  INIT[3941], INIT[3429], INIT[2917], INIT[2405], INIT[1893], INIT[1381], INIT[ 869], INIT[ 357],
  INIT[3940], INIT[3428], INIT[2916], INIT[2404], INIT[1892], INIT[1380], INIT[ 868], INIT[ 356],
  INIT[3939], INIT[3427], INIT[2915], INIT[2403], INIT[1891], INIT[1379], INIT[ 867], INIT[ 355],
  INIT[3938], INIT[3426], INIT[2914], INIT[2402], INIT[1890], INIT[1378], INIT[ 866], INIT[ 354],
  INIT[3937], INIT[3425], INIT[2913], INIT[2401], INIT[1889], INIT[1377], INIT[ 865], INIT[ 353],
  INIT[3936], INIT[3424], INIT[2912], INIT[2400], INIT[1888], INIT[1376], INIT[ 864], INIT[ 352]
};
localparam [255:0] INIT_C = {
  INIT[3999], INIT[3487], INIT[2975], INIT[2463], INIT[1951], INIT[1439], INIT[ 927], INIT[ 415],
  INIT[3998], INIT[3486], INIT[2974], INIT[2462], INIT[1950], INIT[1438], INIT[ 926], INIT[ 414],
  INIT[3997], INIT[3485], INIT[2973], INIT[2461], INIT[1949], INIT[1437], INIT[ 925], INIT[ 413],
  INIT[3996], INIT[3484], INIT[2972], INIT[2460], INIT[1948], INIT[1436], INIT[ 924], INIT[ 412],
  INIT[3995], INIT[3483], INIT[2971], INIT[2459], INIT[1947], INIT[1435], INIT[ 923], INIT[ 411],
  INIT[3994], INIT[3482], INIT[2970], INIT[2458], INIT[1946], INIT[1434], INIT[ 922], INIT[ 410],
  INIT[3993], INIT[3481], INIT[2969], INIT[2457], INIT[1945], INIT[1433], INIT[ 921], INIT[ 409],
  INIT[3992], INIT[3480], INIT[2968], INIT[2456], INIT[1944], INIT[1432], INIT[ 920], INIT[ 408],
  INIT[3991], INIT[3479], INIT[2967], INIT[2455], INIT[1943], INIT[1431], INIT[ 919], INIT[ 407],
  INIT[3990], INIT[3478], INIT[2966], INIT[2454], INIT[1942], INIT[1430], INIT[ 918], INIT[ 406],
  INIT[3989], INIT[3477], INIT[2965], INIT[2453], INIT[1941], INIT[1429], INIT[ 917], INIT[ 405],
  INIT[3988], INIT[3476], INIT[2964], INIT[2452], INIT[1940], INIT[1428], INIT[ 916], INIT[ 404],
  INIT[3987], INIT[3475], INIT[2963], INIT[2451], INIT[1939], INIT[1427], INIT[ 915], INIT[ 403],
  INIT[3986], INIT[3474], INIT[2962], INIT[2450], INIT[1938], INIT[1426], INIT[ 914], INIT[ 402],
  INIT[3985], INIT[3473], INIT[2961], INIT[2449], INIT[1937], INIT[1425], INIT[ 913], INIT[ 401],
  INIT[3984], INIT[3472], INIT[2960], INIT[2448], INIT[1936], INIT[1424], INIT[ 912], INIT[ 400],
  INIT[3983], INIT[3471], INIT[2959], INIT[2447], INIT[1935], INIT[1423], INIT[ 911], INIT[ 399],
  INIT[3982], INIT[3470], INIT[2958], INIT[2446], INIT[1934], INIT[1422], INIT[ 910], INIT[ 398],
  INIT[3981], INIT[3469], INIT[2957], INIT[2445], INIT[1933], INIT[1421], INIT[ 909], INIT[ 397],
  INIT[3980], INIT[3468], INIT[2956], INIT[2444], INIT[1932], INIT[1420], INIT[ 908], INIT[ 396],
  INIT[3979], INIT[3467], INIT[2955], INIT[2443], INIT[1931], INIT[1419], INIT[ 907], INIT[ 395],
  INIT[3978], INIT[3466], INIT[2954], INIT[2442], INIT[1930], INIT[1418], INIT[ 906], INIT[ 394],
  INIT[3977], INIT[3465], INIT[2953], INIT[2441], INIT[1929], INIT[1417], INIT[ 905], INIT[ 393],
  INIT[3976], INIT[3464], INIT[2952], INIT[2440], INIT[1928], INIT[1416], INIT[ 904], INIT[ 392],
  INIT[3975], INIT[3463], INIT[2951], INIT[2439], INIT[1927], INIT[1415], INIT[ 903], INIT[ 391],
  INIT[3974], INIT[3462], INIT[2950], INIT[2438], INIT[1926], INIT[1414], INIT[ 902], INIT[ 390],
  INIT[3973], INIT[3461], INIT[2949], INIT[2437], INIT[1925], INIT[1413], INIT[ 901], INIT[ 389],
  INIT[3972], INIT[3460], INIT[2948], INIT[2436], INIT[1924], INIT[1412], INIT[ 900], INIT[ 388],
  INIT[3971], INIT[3459], INIT[2947], INIT[2435], INIT[1923], INIT[1411], INIT[ 899], INIT[ 387],
  INIT[3970], INIT[3458], INIT[2946], INIT[2434], INIT[1922], INIT[1410], INIT[ 898], INIT[ 386],
  INIT[3969], INIT[3457], INIT[2945], INIT[2433], INIT[1921], INIT[1409], INIT[ 897], INIT[ 385],
  INIT[3968], INIT[3456], INIT[2944], INIT[2432], INIT[1920], INIT[1408], INIT[ 896], INIT[ 384]
};
localparam [255:0] INIT_D = {
  INIT[4031], INIT[3519], INIT[3007], INIT[2495], INIT[1983], INIT[1471], INIT[ 959], INIT[ 447],
  INIT[4030], INIT[3518], INIT[3006], INIT[2494], INIT[1982], INIT[1470], INIT[ 958], INIT[ 446],
  INIT[4029], INIT[3517], INIT[3005], INIT[2493], INIT[1981], INIT[1469], INIT[ 957], INIT[ 445],
  INIT[4028], INIT[3516], INIT[3004], INIT[2492], INIT[1980], INIT[1468], INIT[ 956], INIT[ 444],
  INIT[4027], INIT[3515], INIT[3003], INIT[2491], INIT[1979], INIT[1467], INIT[ 955], INIT[ 443],
  INIT[4026], INIT[3514], INIT[3002], INIT[2490], INIT[1978], INIT[1466], INIT[ 954], INIT[ 442],
  INIT[4025], INIT[3513], INIT[3001], INIT[2489], INIT[1977], INIT[1465], INIT[ 953], INIT[ 441],
  INIT[4024], INIT[3512], INIT[3000], INIT[2488], INIT[1976], INIT[1464], INIT[ 952], INIT[ 440],
  INIT[4023], INIT[3511], INIT[2999], INIT[2487], INIT[1975], INIT[1463], INIT[ 951], INIT[ 439],
  INIT[4022], INIT[3510], INIT[2998], INIT[2486], INIT[1974], INIT[1462], INIT[ 950], INIT[ 438],
  INIT[4021], INIT[3509], INIT[2997], INIT[2485], INIT[1973], INIT[1461], INIT[ 949], INIT[ 437],
  INIT[4020], INIT[3508], INIT[2996], INIT[2484], INIT[1972], INIT[1460], INIT[ 948], INIT[ 436],
  INIT[4019], INIT[3507], INIT[2995], INIT[2483], INIT[1971], INIT[1459], INIT[ 947], INIT[ 435],
  INIT[4018], INIT[3506], INIT[2994], INIT[2482], INIT[1970], INIT[1458], INIT[ 946], INIT[ 434],
  INIT[4017], INIT[3505], INIT[2993], INIT[2481], INIT[1969], INIT[1457], INIT[ 945], INIT[ 433],
  INIT[4016], INIT[3504], INIT[2992], INIT[2480], INIT[1968], INIT[1456], INIT[ 944], INIT[ 432],
  INIT[4015], INIT[3503], INIT[2991], INIT[2479], INIT[1967], INIT[1455], INIT[ 943], INIT[ 431],
  INIT[4014], INIT[3502], INIT[2990], INIT[2478], INIT[1966], INIT[1454], INIT[ 942], INIT[ 430],
  INIT[4013], INIT[3501], INIT[2989], INIT[2477], INIT[1965], INIT[1453], INIT[ 941], INIT[ 429],
  INIT[4012], INIT[3500], INIT[2988], INIT[2476], INIT[1964], INIT[1452], INIT[ 940], INIT[ 428],
  INIT[4011], INIT[3499], INIT[2987], INIT[2475], INIT[1963], INIT[1451], INIT[ 939], INIT[ 427],
  INIT[4010], INIT[3498], INIT[2986], INIT[2474], INIT[1962], INIT[1450], INIT[ 938], INIT[ 426],
  INIT[4009], INIT[3497], INIT[2985], INIT[2473], INIT[1961], INIT[1449], INIT[ 937], INIT[ 425],
  INIT[4008], INIT[3496], INIT[2984], INIT[2472], INIT[1960], INIT[1448], INIT[ 936], INIT[ 424],
  INIT[4007], INIT[3495], INIT[2983], INIT[2471], INIT[1959], INIT[1447], INIT[ 935], INIT[ 423],
  INIT[4006], INIT[3494], INIT[2982], INIT[2470], INIT[1958], INIT[1446], INIT[ 934], INIT[ 422],
  INIT[4005], INIT[3493], INIT[2981], INIT[2469], INIT[1957], INIT[1445], INIT[ 933], INIT[ 421],
  INIT[4004], INIT[3492], INIT[2980], INIT[2468], INIT[1956], INIT[1444], INIT[ 932], INIT[ 420],
  INIT[4003], INIT[3491], INIT[2979], INIT[2467], INIT[1955], INIT[1443], INIT[ 931], INIT[ 419],
  INIT[4002], INIT[3490], INIT[2978], INIT[2466], INIT[1954], INIT[1442], INIT[ 930], INIT[ 418],
  INIT[4001], INIT[3489], INIT[2977], INIT[2465], INIT[1953], INIT[1441], INIT[ 929], INIT[ 417],
  INIT[4000], INIT[3488], INIT[2976], INIT[2464], INIT[1952], INIT[1440], INIT[ 928], INIT[ 416]
};
localparam [255:0] INIT_E = {
  INIT[4063], INIT[3551], INIT[3039], INIT[2527], INIT[2015], INIT[1503], INIT[ 991], INIT[ 479],
  INIT[4062], INIT[3550], INIT[3038], INIT[2526], INIT[2014], INIT[1502], INIT[ 990], INIT[ 478],
  INIT[4061], INIT[3549], INIT[3037], INIT[2525], INIT[2013], INIT[1501], INIT[ 989], INIT[ 477],
  INIT[4060], INIT[3548], INIT[3036], INIT[2524], INIT[2012], INIT[1500], INIT[ 988], INIT[ 476],
  INIT[4059], INIT[3547], INIT[3035], INIT[2523], INIT[2011], INIT[1499], INIT[ 987], INIT[ 475],
  INIT[4058], INIT[3546], INIT[3034], INIT[2522], INIT[2010], INIT[1498], INIT[ 986], INIT[ 474],
  INIT[4057], INIT[3545], INIT[3033], INIT[2521], INIT[2009], INIT[1497], INIT[ 985], INIT[ 473],
  INIT[4056], INIT[3544], INIT[3032], INIT[2520], INIT[2008], INIT[1496], INIT[ 984], INIT[ 472],
  INIT[4055], INIT[3543], INIT[3031], INIT[2519], INIT[2007], INIT[1495], INIT[ 983], INIT[ 471],
  INIT[4054], INIT[3542], INIT[3030], INIT[2518], INIT[2006], INIT[1494], INIT[ 982], INIT[ 470],
  INIT[4053], INIT[3541], INIT[3029], INIT[2517], INIT[2005], INIT[1493], INIT[ 981], INIT[ 469],
  INIT[4052], INIT[3540], INIT[3028], INIT[2516], INIT[2004], INIT[1492], INIT[ 980], INIT[ 468],
  INIT[4051], INIT[3539], INIT[3027], INIT[2515], INIT[2003], INIT[1491], INIT[ 979], INIT[ 467],
  INIT[4050], INIT[3538], INIT[3026], INIT[2514], INIT[2002], INIT[1490], INIT[ 978], INIT[ 466],
  INIT[4049], INIT[3537], INIT[3025], INIT[2513], INIT[2001], INIT[1489], INIT[ 977], INIT[ 465],
  INIT[4048], INIT[3536], INIT[3024], INIT[2512], INIT[2000], INIT[1488], INIT[ 976], INIT[ 464],
  INIT[4047], INIT[3535], INIT[3023], INIT[2511], INIT[1999], INIT[1487], INIT[ 975], INIT[ 463],
  INIT[4046], INIT[3534], INIT[3022], INIT[2510], INIT[1998], INIT[1486], INIT[ 974], INIT[ 462],
  INIT[4045], INIT[3533], INIT[3021], INIT[2509], INIT[1997], INIT[1485], INIT[ 973], INIT[ 461],
  INIT[4044], INIT[3532], INIT[3020], INIT[2508], INIT[1996], INIT[1484], INIT[ 972], INIT[ 460],
  INIT[4043], INIT[3531], INIT[3019], INIT[2507], INIT[1995], INIT[1483], INIT[ 971], INIT[ 459],
  INIT[4042], INIT[3530], INIT[3018], INIT[2506], INIT[1994], INIT[1482], INIT[ 970], INIT[ 458],
  INIT[4041], INIT[3529], INIT[3017], INIT[2505], INIT[1993], INIT[1481], INIT[ 969], INIT[ 457],
  INIT[4040], INIT[3528], INIT[3016], INIT[2504], INIT[1992], INIT[1480], INIT[ 968], INIT[ 456],
  INIT[4039], INIT[3527], INIT[3015], INIT[2503], INIT[1991], INIT[1479], INIT[ 967], INIT[ 455],
  INIT[4038], INIT[3526], INIT[3014], INIT[2502], INIT[1990], INIT[1478], INIT[ 966], INIT[ 454],
  INIT[4037], INIT[3525], INIT[3013], INIT[2501], INIT[1989], INIT[1477], INIT[ 965], INIT[ 453],
  INIT[4036], INIT[3524], INIT[3012], INIT[2500], INIT[1988], INIT[1476], INIT[ 964], INIT[ 452],
  INIT[4035], INIT[3523], INIT[3011], INIT[2499], INIT[1987], INIT[1475], INIT[ 963], INIT[ 451],
  INIT[4034], INIT[3522], INIT[3010], INIT[2498], INIT[1986], INIT[1474], INIT[ 962], INIT[ 450],
  INIT[4033], INIT[3521], INIT[3009], INIT[2497], INIT[1985], INIT[1473], INIT[ 961], INIT[ 449],
  INIT[4032], INIT[3520], INIT[3008], INIT[2496], INIT[1984], INIT[1472], INIT[ 960], INIT[ 448]
};
localparam [255:0] INIT_F = {
  INIT[4095], INIT[3583], INIT[3071], INIT[2559], INIT[2047], INIT[1535], INIT[1023], INIT[ 511],
  INIT[4094], INIT[3582], INIT[3070], INIT[2558], INIT[2046], INIT[1534], INIT[1022], INIT[ 510],
  INIT[4093], INIT[3581], INIT[3069], INIT[2557], INIT[2045], INIT[1533], INIT[1021], INIT[ 509],
  INIT[4092], INIT[3580], INIT[3068], INIT[2556], INIT[2044], INIT[1532], INIT[1020], INIT[ 508],
  INIT[4091], INIT[3579], INIT[3067], INIT[2555], INIT[2043], INIT[1531], INIT[1019], INIT[ 507],
  INIT[4090], INIT[3578], INIT[3066], INIT[2554], INIT[2042], INIT[1530], INIT[1018], INIT[ 506],
  INIT[4089], INIT[3577], INIT[3065], INIT[2553], INIT[2041], INIT[1529], INIT[1017], INIT[ 505],
  INIT[4088], INIT[3576], INIT[3064], INIT[2552], INIT[2040], INIT[1528], INIT[1016], INIT[ 504],
  INIT[4087], INIT[3575], INIT[3063], INIT[2551], INIT[2039], INIT[1527], INIT[1015], INIT[ 503],
  INIT[4086], INIT[3574], INIT[3062], INIT[2550], INIT[2038], INIT[1526], INIT[1014], INIT[ 502],
  INIT[4085], INIT[3573], INIT[3061], INIT[2549], INIT[2037], INIT[1525], INIT[1013], INIT[ 501],
  INIT[4084], INIT[3572], INIT[3060], INIT[2548], INIT[2036], INIT[1524], INIT[1012], INIT[ 500],
  INIT[4083], INIT[3571], INIT[3059], INIT[2547], INIT[2035], INIT[1523], INIT[1011], INIT[ 499],
  INIT[4082], INIT[3570], INIT[3058], INIT[2546], INIT[2034], INIT[1522], INIT[1010], INIT[ 498],
  INIT[4081], INIT[3569], INIT[3057], INIT[2545], INIT[2033], INIT[1521], INIT[1009], INIT[ 497],
  INIT[4080], INIT[3568], INIT[3056], INIT[2544], INIT[2032], INIT[1520], INIT[1008], INIT[ 496],
  INIT[4079], INIT[3567], INIT[3055], INIT[2543], INIT[2031], INIT[1519], INIT[1007], INIT[ 495],
  INIT[4078], INIT[3566], INIT[3054], INIT[2542], INIT[2030], INIT[1518], INIT[1006], INIT[ 494],
  INIT[4077], INIT[3565], INIT[3053], INIT[2541], INIT[2029], INIT[1517], INIT[1005], INIT[ 493],
  INIT[4076], INIT[3564], INIT[3052], INIT[2540], INIT[2028], INIT[1516], INIT[1004], INIT[ 492],
  INIT[4075], INIT[3563], INIT[3051], INIT[2539], INIT[2027], INIT[1515], INIT[1003], INIT[ 491],
  INIT[4074], INIT[3562], INIT[3050], INIT[2538], INIT[2026], INIT[1514], INIT[1002], INIT[ 490],
  INIT[4073], INIT[3561], INIT[3049], INIT[2537], INIT[2025], INIT[1513], INIT[1001], INIT[ 489],
  INIT[4072], INIT[3560], INIT[3048], INIT[2536], INIT[2024], INIT[1512], INIT[1000], INIT[ 488],
  INIT[4071], INIT[3559], INIT[3047], INIT[2535], INIT[2023], INIT[1511], INIT[ 999], INIT[ 487],
  INIT[4070], INIT[3558], INIT[3046], INIT[2534], INIT[2022], INIT[1510], INIT[ 998], INIT[ 486],
  INIT[4069], INIT[3557], INIT[3045], INIT[2533], INIT[2021], INIT[1509], INIT[ 997], INIT[ 485],
  INIT[4068], INIT[3556], INIT[3044], INIT[2532], INIT[2020], INIT[1508], INIT[ 996], INIT[ 484],
  INIT[4067], INIT[3555], INIT[3043], INIT[2531], INIT[2019], INIT[1507], INIT[ 995], INIT[ 483],
  INIT[4066], INIT[3554], INIT[3042], INIT[2530], INIT[2018], INIT[1506], INIT[ 994], INIT[ 482],
  INIT[4065], INIT[3553], INIT[3041], INIT[2529], INIT[2017], INIT[1505], INIT[ 993], INIT[ 481],
  INIT[4064], INIT[3552], INIT[3040], INIT[2528], INIT[2016], INIT[1504], INIT[ 992], INIT[ 480]
};
